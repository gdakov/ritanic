/*
Copyright 2022-2024 Goran Dakov, D.O.B. 11 January 1983, lives in Bristol UK in 2024

Licensed under GPL v3 or commercial license.

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/


(* align_width=C,A_out/2,B_out/2 align_height=R *) module fpucadd_compress_24(clk,R,C,A_out,B_out);
  input pwire clk;
  input pwire [23:0] R;
  input pwire [23:0] C;
  output pwire [47:0] A_out;
  output pwire [47:0] B_out;
  (* register *) reg REGS_0;
  (* register *) reg REGS_1;
  (* register *) reg REGS_2;
  (* register *) reg REGS_3;
  (* register *) reg REGS_4;
  (* register *) reg REGS_5;
  (* register *) reg REGS_6;
  (* register *) reg REGS_7;
  (* register *) reg REGS_8;
  (* register *) reg REGS_9;
  (* register *) reg REGS_10;
  (* register *) reg REGS_11;
  (* register *) reg REGS_12;
  (* register *) reg REGS_13;
  (* register *) reg REGS_14;
  (* register *) reg REGS_15;
  (* register *) reg REGS_16;
  (* register *) reg REGS_17;
  (* register *) reg REGS_18;
  (* register *) reg REGS_19;
  (* register *) reg REGS_20;
  (* register *) reg REGS_21;
  (* register *) reg REGS_22;
  (* register *) reg REGS_23;
  (* register *) reg REGS_24;
  (* register *) reg REGS_25;
  (* register *) reg REGS_26;
  (* register *) reg REGS_27;
  (* register *) reg REGS_28;
  (* register *) reg REGS_29;
  (* register *) reg REGS_30;
  (* register *) reg REGS_31;
  (* register *) reg REGS_32;
  (* register *) reg REGS_33;
  (* register *) reg REGS_34;
  (* register *) reg REGS_35;
  (* register *) reg REGS_36;
  (* register *) reg REGS_37;
  (* register *) reg REGS_38;
  (* register *) reg REGS_39;
  (* register *) reg REGS_40;
  (* register *) reg REGS_41;
  (* register *) reg REGS_42;
  (* register *) reg REGS_43;
  (* register *) reg REGS_44;
  (* register *) reg REGS_45;
  (* register *) reg REGS_46;
  (* register *) reg REGS_47;
  (* register *) reg REGS_48;
  (* register *) reg REGS_49;
  (* register *) reg REGS_50;
  (* register *) reg REGS_51;
  (* register *) reg REGS_52;
  (* register *) reg REGS_53;
  (* register *) reg REGS_54;
  (* register *) reg REGS_55;
  (* register *) reg REGS_56;
  (* register *) reg REGS_57;
  (* register *) reg REGS_58;
  (* register *) reg REGS_59;
  (* register *) reg REGS_60;
  (* register *) reg REGS_61;
  (* register *) reg REGS_62;
  (* register *) reg REGS_63;
  (* register *) reg REGS_64;
  (* register *) reg REGS_65;
  (* register *) reg REGS_66;
  (* register *) reg REGS_67;
  (* register *) reg REGS_68;
  (* register *) reg REGS_69;
  (* register *) reg REGS_70;
  (* register *) reg REGS_71;
  (* register *) reg REGS_72;
  (* register *) reg REGS_73;
  (* register *) reg REGS_74;
  (* register *) reg REGS_75;
  (* register *) reg REGS_76;
  (* register *) reg REGS_77;
  (* register *) reg REGS_78;
  (* register *) reg REGS_79;
  (* register *) reg REGS_80;
  (* register *) reg REGS_81;
  (* register *) reg REGS_82;
  (* register *) reg REGS_83;
  (* register *) reg REGS_84;
  (* register *) reg REGS_85;
  (* register *) reg REGS_86;
  (* register *) reg REGS_87;
  (* register *) reg REGS_88;
  (* register *) reg REGS_89;
  (* register *) reg REGS_90;
  (* register *) reg REGS_91;
  (* register *) reg REGS_92;
  (* register *) reg REGS_93;
  (* register *) reg REGS_94;
  (* register *) reg REGS_95;
  (* register *) reg REGS_96;
  (* register *) reg REGS_97;
  (* register *) reg REGS_98;
  (* register *) reg REGS_99;
  (* register *) reg REGS_100;
  (* register *) reg REGS_101;
  (* register *) reg REGS_102;
  (* register *) reg REGS_103;
  (* register *) reg REGS_104;
  (* register *) reg REGS_105;
  (* register *) reg REGS_106;
  (* register *) reg REGS_107;
  (* register *) reg REGS_108;
  (* register *) reg REGS_109;
  (* register *) reg REGS_110;
  (* register *) reg REGS_111;
  (* register *) reg REGS_112;
  (* register *) reg REGS_113;
  (* register *) reg REGS_114;
  (* register *) reg REGS_115;
  (* register *) reg REGS_116;
  (* register *) reg REGS_117;
  (* register *) reg REGS_118;
  (* register *) reg REGS_119;
  (* register *) reg REGS_120;
  (* register *) reg REGS_121;
  (* register *) reg REGS_122;
  (* register *) reg REGS_123;
  (* register *) reg REGS_124;
  (* register *) reg REGS_125;
  (* register *) reg REGS_126;
  (* register *) reg REGS_127;
  (* register *) reg REGS_128;
  (* register *) reg REGS_129;
  (* register *) reg REGS_130;
  (* register *) reg REGS_131;
  (* register *) reg REGS_132;
  (* register *) reg REGS_133;
  (* register *) reg REGS_134;
  (* register *) reg REGS_135;
  (* register *) reg REGS_136;
  (* register *) reg REGS_137;
  (* register *) reg REGS_138;
  (* register *) reg REGS_139;
  (* register *) reg REGS_140;
  (* register *) reg REGS_141;
  (* register *) reg REGS_142;
  (* register *) reg REGS_143;
  (* register *) reg REGS_144;
  (* register *) reg REGS_145;
  (* register *) reg REGS_146;
  (* register *) reg REGS_147;
  (* register *) reg REGS_148;
  (* register *) reg REGS_149;
  (* register *) reg REGS_150;
  (* register *) reg REGS_151;
  (* register *) reg REGS_152;
  (* register *) reg REGS_153;
  (* register *) reg REGS_154;
  (* register *) reg REGS_155;
  (* register *) reg REGS_156;
  (* register *) reg REGS_157;
  (* register *) reg REGS_158;
  (* register *) reg REGS_159;
  (* register *) reg REGS_160;
  (* register *) reg REGS_161;
  (* register *) reg REGS_162;
  (* register *) reg REGS_163;
  (* register *) reg REGS_164;
  (* register *) reg REGS_165;
  (* register *) reg REGS_166;
  (* register *) reg REGS_167;
  (* register *) reg REGS_168;
  (* register *) reg REGS_169;
  (* register *) reg REGS_170;
  (* register *) reg REGS_171;
  (* register *) reg REGS_172;
  (* register *) reg REGS_173;
  (* register *) reg REGS_174;
  (* register *) reg REGS_175;
  (* register *) reg REGS_176;
  (* register *) reg REGS_177;
  (* register *) reg REGS_178;
  (* register *) reg REGS_179;
  (* register *) reg REGS_180;
  (* register *) reg REGS_181;
  (* register *) reg REGS_182;
  (* register *) reg REGS_183;
  (* register *) reg REGS_184;
  (* register *) reg REGS_185;
  (* register *) reg REGS_186;
  (* register *) reg REGS_187;
  (* register *) reg REGS_188;
  (* register *) reg REGS_189;
  (* register *) reg REGS_190;
  (* register *) reg REGS_191;
  (* register *) reg REGS_192;
  (* register *) reg REGS_193;
  (* register *) reg REGS_194;
  (* register *) reg REGS_195;
  (* register *) reg REGS_196;
  (* register *) reg REGS_197;
  (* register *) reg REGS_198;
  (* register *) reg REGS_199;
  (* register *) reg REGS_200;
  (* register *) reg REGS_201;
  (* register *) reg REGS_202;
  (* register *) reg REGS_203;
  (* register *) reg REGS_204;
  (* register *) reg REGS_205;
  (* register *) reg REGS_206;
  (* register *) reg REGS_207;
  (* register *) reg REGS_208;
  (* register *) reg REGS_209;
  (* register *) reg REGS_210;
  (* register *) reg REGS_211;
  (* register *) reg REGS_212;
  (* register *) reg REGS_213;
  (* register *) reg REGS_214;
  (* register *) reg REGS_215;
  (* register *) reg REGS_216;
  (* register *) reg REGS_217;
  (* register *) reg REGS_218;
  (* register *) reg REGS_219;
  (* register *) reg REGS_220;
  (* register *) reg REGS_221;
  (* register *) reg REGS_222;
  (* register *) reg REGS_223;
  (* register *) reg REGS_224;
  (* register *) reg REGS_225;
  (* register *) reg REGS_226;
  (* register *) reg REGS_227;
  (* register *) reg REGS_228;
  (* register *) reg REGS_229;
  (* register *) reg REGS_230;
  (* register *) reg REGS_231;
  (* register *) reg REGS_232;
  (* register *) reg REGS_233;
  (* register *) reg REGS_234;
  (* register *) reg REGS_235;
  (* register *) reg REGS_236;
  (* register *) reg REGS_237;
  (* register *) reg REGS_238;
  (* register *) reg REGS_239;
  (* register *) reg REGS_240;
  (* register *) reg REGS_241;
  (* register *) reg REGS_242;
  (* register *) reg REGS_243;
  (* register *) reg REGS_244;
  (* register *) reg REGS_245;
  (* register *) reg REGS_246;
  (* register *) reg REGS_247;
  (* register *) reg REGS_248;
  (* register *) reg REGS_249;
  (* register *) reg REGS_250;
  (* register *) reg REGS_251;
  (* register *) reg REGS_252;
  (* register *) reg REGS_253;
  (* register *) reg REGS_254;
  (* register *) reg REGS_255;
  (* register *) reg REGS_256;
  (* register *) reg REGS_257;
  (* register *) reg REGS_258;
  (* register *) reg REGS_259;
  (* register *) reg REGS_260;
  (* register *) reg REGS_261;
  (* register *) reg REGS_262;
  (* register *) reg REGS_263;
  (* register *) reg REGS_264;
  (* register *) reg REGS_265;
  (* register *) reg REGS_266;
  (* register *) reg REGS_267;
  (* register *) reg REGS_268;
  (* register *) reg REGS_269;
  (* register *) reg REGS_270;
  (* register *) reg REGS_271;
  (* register *) reg REGS_272;
  (* register *) reg REGS_273;
  (* register *) reg REGS_274;
  (* register *) reg REGS_275;
  (* register *) reg REGS_276;
  (* register *) reg REGS_277;
  (* register *) reg REGS_278;
  (* register *) reg REGS_279;
  (* register *) reg REGS_280;
  (* register *) reg REGS_281;
  (* register *) reg REGS_282;
  (* register *) reg REGS_283;
  (* register *) reg REGS_284;
  (* register *) reg REGS_285;
  (* register *) reg REGS_286;
  (* register *) reg REGS_287;
  (* register *) reg REGS_288;
  (* register *) reg REGS_289;
  (* register *) reg REGS_290;
  (* register *) reg REGS_291;
  (* register *) reg REGS_292;
  (* register *) reg REGS_293;
  (* register *) reg REGS_294;
  (* register *) reg REGS_295;
  (* register *) reg REGS_296;
  (* register *) reg REGS_297;
  (* register *) reg REGS_298;
  (* register *) reg REGS_299;
  (* register *) reg REGS_300;
  (* register *) reg REGS_301;
  (* register *) reg REGS_302;
  (* register *) reg REGS_303;
  (* register *) reg REGS_304;
  (* register *) reg REGS_305;
  (* register *) reg REGS_306;
  (* register *) reg REGS_307;
  (* register *) reg REGS_308;
  (* register *) reg REGS_309;
  (* register *) reg REGS_310;
  (* register *) reg REGS_311;
  (* register *) reg REGS_312;
  (* register *) reg REGS_313;
  (* register *) reg REGS_314;
  (* register *) reg REGS_315;
  (* register *) reg REGS_316;
  (* register *) reg REGS_317;
  (* register *) reg REGS_318;
  (* register *) reg REGS_319;
  (* register *) reg REGS_320;
  (* register *) reg REGS_321;
  (* register *) reg REGS_322;
  (* register *) reg REGS_323;
  (* register *) reg REGS_324;
  (* register *) reg REGS_325;
  (* register *) reg REGS_326;
  (* register *) reg REGS_327;
  (* register *) reg REGS_328;
  (* register *) reg REGS_329;
  (* register *) reg REGS_330;
  (* register *) reg REGS_331;
  (* register *) reg REGS_332;
  (* register *) reg REGS_333;
  (* register *) reg REGS_334;
  (* register *) reg REGS_335;
  (* register *) reg REGS_336;
  (* register *) reg REGS_337;
  (* register *) reg REGS_338;
  (* register *) reg REGS_339;
  (* register *) reg REGS_340;
  (* register *) reg REGS_341;
  (* register *) reg REGS_342;
  (* register *) reg REGS_343;
  (* register *) reg REGS_344;
  (* register *) reg REGS_345;
  (* register *) reg REGS_346;
  (* register *) reg REGS_347;
  (* register *) reg REGS_348;
  (* register *) reg REGS_349;
  (* register *) reg REGS_350;
  (* register *) reg REGS_351;
  (* register *) reg REGS_352;
  (* register *) reg REGS_353;
  (* register *) reg REGS_354;
  (* register *) reg REGS_355;
  (* register *) reg REGS_356;
  (* register *) reg REGS_357;
  (* register *) reg REGS_358;
  (* register *) reg REGS_359;
  (* register *) reg REGS_360;
  (* register *) reg REGS_361;
  (* register *) reg REGS_362;
  (* register *) reg REGS_363;
  (* register *) reg REGS_364;
  (* register *) reg REGS_365;
  (* register *) reg REGS_366;
  (* register *) reg REGS_367;
  (* register *) reg REGS_368;
  (* register *) reg REGS_369;
  (* register *) reg REGS_370;
  (* register *) reg REGS_371;
  (* register *) reg REGS_372;
  (* register *) reg REGS_373;
  (* register *) reg REGS_374;
  (* register *) reg REGS_375;
  (* register *) reg REGS_376;
  (* register *) reg REGS_377;
  (* register *) reg REGS_378;
  (* register *) reg REGS_379;
  (* register *) reg REGS_380;
  (* register *) reg REGS_381;
  (* register *) reg REGS_382;
  (* register *) pwire FA_out_0;
  (* register *) pwire FA_out_1;
  (* register *) pwire FA_out_2;
  (* register *) pwire FA_out_3;
  (* register *) pwire FA_out_4;
  (* register *) pwire FA_out_5;
  (* register *) pwire FA_out_6;
  (* register *) pwire FA_out_7;
  (* register *) pwire FA_out_8;
  (* register *) pwire FA_out_9;
  (* register *) pwire FA_out_10;
  (* register *) pwire FA_out_11;
  (* register *) pwire FA_out_12;
  (* register *) pwire FA_out_13;
  (* register *) pwire FA_out_14;
  (* register *) pwire FA_out_15;
  (* register *) pwire FA_out_16;
  (* register *) pwire FA_out_17;
  (* register *) pwire FA_out_18;
  (* register *) pwire FA_out_19;
  (* register *) pwire FA_out_20;
  (* register *) pwire FA_out_21;
  (* register *) pwire FA_out_22;
  (* register *) pwire FA_out_23;
  (* register *) pwire FA_out_24;
  (* register *) pwire FA_out_25;
  (* register *) pwire FA_out_26;
  (* register *) pwire FA_out_27;
  (* register *) pwire FA_out_28;
  (* register *) pwire FA_out_29;
  (* register *) pwire FA_out_30;
  (* register *) pwire FA_out_31;
  (* register *) pwire FA_out_32;
  (* register *) pwire FA_out_33;
  (* register *) pwire FA_out_34;
  (* register *) pwire FA_out_35;
  (* register *) pwire FA_out_36;
  (* register *) pwire FA_out_37;
  (* register *) pwire FA_out_38;
  (* register *) pwire FA_out_39;
  (* register *) pwire FA_out_40;
  (* register *) pwire FA_out_41;
  (* register *) pwire FA_out_42;
  (* register *) pwire FA_out_43;
  (* register *) pwire FA_out_44;
  (* register *) pwire FA_out_45;
  (* register *) pwire FA_out_46;
  (* register *) pwire FA_out_47;
  (* register *) pwire FA_out_48;
  (* register *) pwire FA_out_49;
  (* register *) pwire FA_out_50;
  (* register *) pwire FA_out_51;
  (* register *) pwire FA_out_52;
  (* register *) pwire FA_out_53;
  (* register *) pwire FA_out_54;
  (* register *) pwire FA_out_55;
  (* register *) pwire FA_out_56;
  (* register *) pwire FA_out_57;
  (* register *) pwire FA_out_58;
  (* register *) pwire FA_out_59;
  (* register *) pwire FA_out_60;
  (* register *) pwire FA_out_61;
  (* register *) pwire FA_out_62;
  (* register *) pwire FA_out_63;
  (* register *) pwire FA_out_64;
  (* register *) pwire FA_out_65;
  (* register *) pwire FA_out_66;
  (* register *) pwire FA_out_67;
  (* register *) pwire FA_out_68;
  (* register *) pwire FA_out_69;
  (* register *) pwire FA_out_70;
  (* register *) pwire FA_out_71;
  (* register *) pwire FA_out_72;
  (* register *) pwire FA_out_73;
  (* register *) pwire FA_out_74;
  (* register *) pwire FA_out_75;
  (* register *) pwire FA_out_76;
  (* register *) pwire FA_out_77;
  (* register *) pwire FA_out_78;
  (* register *) pwire FA_out_79;
  (* register *) pwire FA_out_80;
  (* register *) pwire FA_out_81;
  (* register *) pwire FA_out_82;
  (* register *) pwire FA_out_83;
  (* register *) pwire FA_out_84;
  (* register *) pwire FA_out_85;
  (* register *) pwire FA_out_86;
  (* register *) pwire FA_out_87;
  (* register *) pwire FA_out_88;
  (* register *) pwire FA_out_89;
  (* register *) pwire FA_out_90;
  (* register *) pwire FA_out_91;
  (* register *) pwire FA_out_92;
  (* register *) pwire FA_out_93;
  (* register *) pwire FA_out_94;
  (* register *) pwire FA_out_95;
  (* register *) pwire FA_out_96;
  (* register *) pwire FA_out_97;
  (* register *) pwire FA_out_98;
  (* register *) pwire FA_out_99;
  (* register *) pwire FA_out_100;
  (* register *) pwire FA_out_101;
  (* register *) pwire FA_out_102;
  (* register *) pwire FA_out_103;
  (* register *) pwire FA_out_104;
  (* register *) pwire FA_out_105;
  (* register *) pwire FA_out_106;
  (* register *) pwire FA_out_107;
  (* register *) pwire FA_out_108;
  (* register *) pwire FA_out_109;
  (* register *) pwire FA_out_110;
  (* register *) pwire FA_out_111;
  (* register *) pwire FA_out_112;
  (* register *) pwire FA_out_113;
  (* register *) pwire FA_out_114;
  (* register *) pwire FA_out_115;
  (* register *) pwire FA_out_116;
  (* register *) pwire FA_out_117;
  (* register *) pwire FA_out_118;
  (* register *) pwire FA_out_119;
  (* register *) pwire FA_out_120;
  (* register *) pwire FA_out_121;
  (* register *) pwire FA_out_122;
  (* register *) pwire FA_out_123;
  (* register *) pwire FA_out_124;
  (* register *) pwire FA_out_125;
  (* register *) pwire FA_out_126;
  (* register *) pwire FA_out_127;
  (* register *) pwire FA_out_128;
  (* register *) pwire FA_out_129;
  (* register *) pwire FA_out_130;
  (* register *) pwire FA_out_131;
  (* register *) pwire FA_out_132;
  (* register *) pwire FA_out_133;
  (* register *) pwire FA_out_134;
  (* register *) pwire FA_out_135;
  (* register *) pwire FA_out_136;
  (* register *) pwire FA_out_137;
  (* register *) pwire FA_out_138;
  (* register *) pwire FA_out_139;
  (* register *) pwire FA_out_140;
  (* register *) pwire FA_out_141;
  (* register *) pwire FA_out_142;
  (* register *) pwire FA_out_143;
  (* register *) pwire FA_out_144;
  (* register *) pwire FA_out_145;
  (* register *) pwire FA_out_146;
  (* register *) pwire FA_out_147;
  (* register *) pwire FA_out_148;
  (* register *) pwire FA_out_149;
  (* register *) pwire FA_out_150;
  (* register *) pwire FA_out_151;
  (* register *) pwire FA_out_152;
  (* register *) pwire FA_out_153;
  (* register *) pwire FA_out_154;
  (* register *) pwire FA_out_155;
  (* register *) pwire FA_out_156;
  (* register *) pwire FA_out_157;
  (* register *) pwire FA_out_158;
  (* register *) pwire FA_out_159;
  (* register *) pwire FA_out_160;
  (* register *) pwire FA_out_161;
  (* register *) pwire FA_out_162;
  (* register *) pwire FA_out_163;
  (* register *) pwire FA_out_164;
  (* register *) pwire FA_out_165;
  (* register *) pwire FA_out_166;
  (* register *) pwire FA_out_167;
  (* register *) pwire FA_out_168;
  (* register *) pwire FA_out_169;
  (* register *) pwire FA_out_170;
  (* register *) pwire FA_out_171;
  (* register *) pwire FA_out_172;
  (* register *) pwire FA_out_173;
  (* register *) pwire FA_out_174;
  (* register *) pwire FA_out_175;
  (* register *) pwire FA_out_176;
  (* register *) pwire FA_out_177;
  (* register *) pwire FA_out_178;
  (* register *) pwire FA_out_179;
  (* register *) pwire FA_out_180;
  (* register *) pwire FA_out_181;
  (* register *) pwire FA_out_182;
  (* register *) pwire FA_out_183;
  (* register *) pwire FA_out_184;
  (* register *) pwire FA_out_185;
  (* register *) pwire FA_out_186;
  (* register *) pwire FA_out_187;
  (* register *) pwire FA_out_188;
  (* register *) pwire FA_out_189;
  (* register *) pwire FA_out_190;
  (* register *) pwire FA_out_191;
  (* register *) pwire FA_out_192;
  (* register *) pwire FA_out_193;
  (* register *) pwire FA_out_194;
  (* register *) pwire FA_out_195;
  (* register *) pwire FA_out_196;
  (* register *) pwire FA_out_197;
  (* register *) pwire FA_out_198;
  (* register *) pwire FA_out_199;
  (* register *) pwire FA_out_200;
  (* register *) pwire FA_out_201;
  (* register *) pwire FA_out_202;
  (* register *) pwire FA_out_203;
  (* register *) pwire FA_out_204;
  (* register *) pwire FA_out_205;
  (* register *) pwire FA_out_206;
  (* register *) pwire FA_out_207;
  (* register *) pwire FA_out_208;
  (* register *) pwire FA_out_209;
  (* register *) pwire FA_out_210;
  (* register *) pwire FA_out_211;
  (* register *) pwire FA_out_212;
  (* register *) pwire FA_out_213;
  (* register *) pwire FA_out_214;
  (* register *) pwire FA_out_215;
  (* register *) pwire FA_out_216;
  (* register *) pwire FA_out_217;
  (* register *) pwire FA_out_218;
  (* register *) pwire FA_out_219;
  (* register *) pwire FA_out_220;
  (* register *) pwire FA_out_221;
  (* register *) pwire FA_out_222;
  (* register *) pwire FA_out_223;
  (* register *) pwire FA_out_224;
  (* register *) pwire FA_out_225;
  (* register *) pwire FA_out_226;
  (* register *) pwire FA_out_227;
  (* register *) pwire FA_out_228;
  (* register *) pwire FA_out_229;
  (* register *) pwire FA_out_230;
  (* register *) pwire FA_out_231;
  (* register *) pwire FA_out_232;
  (* register *) pwire FA_out_233;
  (* register *) pwire FA_out_234;
  (* register *) pwire FA_out_235;
  (* register *) pwire FA_out_236;
  (* register *) pwire FA_out_237;
  (* register *) pwire FA_out_238;
  (* register *) pwire FA_out_239;
  (* register *) pwire FA_out_240;
  (* register *) pwire FA_out_241;
  (* register *) pwire FA_out_242;
  (* register *) pwire FA_out_243;
  (* register *) pwire FA_out_244;
  (* register *) pwire FA_out_245;
  (* register *) pwire FA_out_246;
  (* register *) pwire FA_out_247;
  (* register *) pwire FA_out_248;
  (* register *) pwire FA_out_249;
  (* register *) pwire FA_out_250;
  (* register *) pwire FA_out_251;
  (* register *) pwire FA_out_252;
  (* register *) pwire FA_out_253;
  (* register *) pwire FA_out_254;
  (* register *) pwire FA_out_255;
  (* register *) pwire FA_out_256;
  (* register *) pwire FA_out_257;
  (* register *) pwire FA_out_258;
  (* register *) pwire FA_out_259;
  (* register *) pwire FA_out_260;
  (* register *) pwire FA_out_261;
  (* register *) pwire FA_out_262;
  (* register *) pwire FA_out_263;
  (* register *) pwire FA_out_264;
  (* register *) pwire FA_out_265;
  (* register *) pwire FA_out_266;
  (* register *) pwire FA_out_267;
  (* register *) pwire FA_out_268;
  (* register *) pwire FA_out_269;
  (* register *) pwire FA_out_270;
  (* register *) pwire FA_out_271;
  (* register *) pwire FA_out_272;
  (* register *) pwire FA_out_273;
  (* register *) pwire FA_out_274;
  (* register *) pwire FA_out_275;
  (* register *) pwire FA_out_276;
  (* register *) pwire FA_out_277;
  (* register *) pwire FA_out_278;
  (* register *) pwire FA_out_279;
  (* register *) pwire FA_out_280;
  (* register *) pwire FA_out_281;
  (* register *) pwire FA_out_282;
  (* register *) pwire FA_out_283;
  (* register *) pwire FA_out_284;
  (* register *) pwire FA_out_285;
  (* register *) pwire FA_out_286;
  (* register *) pwire FA_out_287;
  (* register *) pwire FA_out_288;
  (* register *) pwire FA_out_289;
  (* register *) pwire FA_out_290;
  (* register *) pwire FA_out_291;
  (* register *) pwire FA_out_292;
  (* register *) pwire FA_out_293;
  (* register *) pwire FA_out_294;
  (* register *) pwire FA_out_295;
  (* register *) pwire FA_out_296;
  (* register *) pwire FA_out_297;
  (* register *) pwire FA_out_298;
  (* register *) pwire FA_out_299;
  (* register *) pwire FA_out_300;
  (* register *) pwire FA_out_301;
  (* register *) pwire FA_out_302;
  (* register *) pwire FA_out_303;
  (* register *) pwire FA_out_304;
  (* register *) pwire FA_out_305;
  (* register *) pwire FA_out_306;
  (* register *) pwire FA_out_307;
  (* register *) pwire FA_out_308;
  (* register *) pwire FA_out_309;
  (* register *) pwire FA_out_310;
  (* register *) pwire FA_out_311;
  (* register *) pwire FA_out_312;
  (* register *) pwire FA_out_313;
  (* register *) pwire FA_out_314;
  (* register *) pwire FA_out_315;
  (* register *) pwire FA_out_316;
  (* register *) pwire FA_out_317;
  (* register *) pwire FA_out_318;
  (* register *) pwire FA_out_319;
  (* register *) pwire FA_out_320;
  (* register *) pwire FA_out_321;
  (* register *) pwire FA_out_322;
  (* register *) pwire FA_out_323;
  (* register *) pwire FA_out_324;
  (* register *) pwire FA_out_325;
  (* register *) pwire FA_out_326;
  (* register *) pwire FA_out_327;
  (* register *) pwire FA_out_328;
  (* register *) pwire FA_out_329;
  (* register *) pwire FA_out_330;
  (* register *) pwire FA_out_331;
  (* register *) pwire FA_out_332;
  (* register *) pwire FA_out_333;
  (* register *) pwire FA_out_334;
  (* register *) pwire FA_out_335;
  (* register *) pwire FA_out_336;
  (* register *) pwire FA_out_337;
  (* register *) pwire FA_out_338;
  (* register *) pwire FA_out_339;
  (* register *) pwire FA_out_340;
  (* register *) pwire FA_out_341;
  (* register *) pwire FA_out_342;
  (* register *) pwire FA_out_343;
  (* register *) pwire FA_out_344;
  (* register *) pwire FA_out_345;
  (* register *) pwire FA_out_346;
  (* register *) pwire FA_out_347;
  (* register *) pwire FA_out_348;
  (* register *) pwire FA_out_349;
  (* register *) pwire FA_out_350;
  (* register *) pwire FA_out_351;
  (* register *) pwire FA_out_352;
  (* register *) pwire FA_out_353;
  (* register *) pwire FA_out_354;
  (* register *) pwire FA_out_355;
  (* register *) pwire FA_out_356;
  (* register *) pwire FA_out_357;
  (* register *) pwire FA_out_358;
  (* register *) pwire FA_out_359;
  (* register *) pwire FA_out_360;
  (* register *) pwire FA_out_361;
  (* register *) pwire FA_out_362;
  (* register *) pwire FA_out_363;
  (* register *) pwire FA_out_364;
  (* register *) pwire FA_out_365;
  (* register *) pwire FA_out_366;
  (* register *) pwire FA_out_367;
  (* register *) pwire FA_out_368;
  (* register *) pwire FA_out_369;
  (* register *) pwire FA_out_370;
  (* register *) pwire FA_out_371;
  (* register *) pwire FA_out_372;
  (* register *) pwire FA_out_373;
  (* register *) pwire FA_out_374;
  (* register *) pwire FA_out_375;
  (* register *) pwire FA_out_376;
  (* register *) pwire FA_out_377;
  (* register *) pwire FA_out_378;
  (* register *) pwire FA_out_379;
  (* register *) pwire FA_out_380;
  (* register *) pwire FA_out_381;
  (* register *) pwire FA_out_382;
  (* register *) pwire FA_out_383;
  (* register *) pwire FA_out_384;
  (* register *) pwire FA_out_385;
  (* register *) pwire FA_out_386;
  (* register *) pwire FA_out_387;
  (* register *) pwire FA_out_388;
  (* register *) pwire FA_out_389;
  (* register *) pwire FA_out_390;
  (* register *) pwire FA_out_391;
  (* register *) pwire FA_out_392;
  (* register *) pwire FA_out_393;
  (* register *) pwire FA_out_394;
  (* register *) pwire FA_out_395;
  (* register *) pwire FA_out_396;
  (* register *) pwire FA_out_397;
  (* register *) pwire FA_out_398;
  (* register *) pwire FA_out_399;
  (* register *) pwire FA_out_400;
  (* register *) pwire FA_out_401;
  (* register *) pwire FA_out_402;
  (* register *) pwire FA_out_403;
  (* register *) pwire FA_out_404;
  (* register *) pwire FA_out_405;
  (* register *) pwire FA_out_406;
  (* register *) pwire FA_out_407;
  (* register *) pwire FA_out_408;
  (* register *) pwire FA_out_409;
  (* register *) pwire FA_out_410;
  (* register *) pwire FA_out_411;
  (* register *) pwire FA_out_412;
  (* register *) pwire FA_out_413;
  (* register *) pwire FA_out_414;
  (* register *) pwire FA_out_415;
  (* register *) pwire FA_out_416;
  (* register *) pwire FA_out_417;
  (* register *) pwire FA_out_418;
  (* register *) pwire FA_out_419;
  (* register *) pwire FA_out_420;
  (* register *) pwire FA_out_421;
  (* register *) pwire FA_out_422;
  (* register *) pwire FA_out_423;
  (* register *) pwire FA_out_424;
  (* register *) pwire FA_out_425;
  (* register *) pwire FA_out_426;
  (* register *) pwire FA_out_427;
  (* register *) pwire FA_out_428;
  (* register *) pwire FA_out_429;
  (* register *) pwire FA_out_430;
  (* register *) pwire FA_out_431;
  (* register *) pwire FA_out_432;
  (* register *) pwire FA_out_433;
  (* register *) pwire FA_out_434;
  (* register *) pwire FA_out_435;
  (* register *) pwire FA_out_436;
  (* register *) pwire FA_out_437;
  (* register *) pwire FA_out_438;
  (* register *) pwire FA_out_439;
  (* register *) pwire FA_out_440;
  (* register *) pwire FA_out_441;
  (* register *) pwire FA_out_442;
  (* register *) pwire FA_out_443;
  (* register *) pwire FA_out_444;
  (* register *) pwire FA_out_445;
  (* register *) pwire FA_out_446;
  (* register *) pwire FA_out_447;
  (* register *) pwire FA_out_448;
  (* register *) pwire FA_out_449;
  (* register *) pwire FA_out_450;
  (* register *) pwire FA_out_451;
  (* register *) pwire FA_out_452;
  (* register *) pwire FA_out_453;
  (* register *) pwire FA_out_454;
  (* register *) pwire FA_out_455;
  (* register *) pwire FA_out_456;
  (* register *) pwire FA_out_457;
  (* register *) pwire FA_out_458;
  (* register *) pwire FA_out_459;
  (* register *) pwire FA_out_460;
  (* register *) pwire FA_out_461;
  (* register *) pwire FA_out_462;
  (* register *) pwire FA_out_463;
  (* register *) pwire FA_out_464;
  (* register *) pwire FA_out_465;
  (* register *) pwire FA_out_466;
  (* register *) pwire FA_out_467;
  (* register *) pwire FA_out_468;
  (* register *) pwire FA_out_469;
  (* register *) pwire FA_out_470;
  (* register *) pwire FA_out_471;
  (* register *) pwire FA_out_472;
  (* register *) pwire FA_out_473;
  (* register *) pwire FA_out_474;
  (* register *) pwire FA_out_475;
  (* register *) pwire FA_out_476;
  (* register *) pwire FA_out_477;
  (* register *) pwire FA_out_478;
  (* register *) pwire FA_out_479;
  (* register *) pwire FA_out_480;
  (* register *) pwire FA_out_481;
  (* register *) pwire FA_out_482;
  (* register *) pwire FA_out_483;
  (* register *) pwire FA_cout_0;
  (* register *) pwire FA_cout_1;
  (* register *) pwire FA_cout_2;
  (* register *) pwire FA_cout_3;
  (* register *) pwire FA_cout_4;
  (* register *) pwire FA_cout_5;
  (* register *) pwire FA_cout_6;
  (* register *) pwire FA_cout_7;
  (* register *) pwire FA_cout_8;
  (* register *) pwire FA_cout_9;
  (* register *) pwire FA_cout_10;
  (* register *) pwire FA_cout_11;
  (* register *) pwire FA_cout_12;
  (* register *) pwire FA_cout_13;
  (* register *) pwire FA_cout_14;
  (* register *) pwire FA_cout_15;
  (* register *) pwire FA_cout_16;
  (* register *) pwire FA_cout_17;
  (* register *) pwire FA_cout_18;
  (* register *) pwire FA_cout_19;
  (* register *) pwire FA_cout_20;
  (* register *) pwire FA_cout_21;
  (* register *) pwire FA_cout_22;
  (* register *) pwire FA_cout_23;
  (* register *) pwire FA_cout_24;
  (* register *) pwire FA_cout_25;
  (* register *) pwire FA_cout_26;
  (* register *) pwire FA_cout_27;
  (* register *) pwire FA_cout_28;
  (* register *) pwire FA_cout_29;
  (* register *) pwire FA_cout_30;
  (* register *) pwire FA_cout_31;
  (* register *) pwire FA_cout_32;
  (* register *) pwire FA_cout_33;
  (* register *) pwire FA_cout_34;
  (* register *) pwire FA_cout_35;
  (* register *) pwire FA_cout_36;
  (* register *) pwire FA_cout_37;
  (* register *) pwire FA_cout_38;
  (* register *) pwire FA_cout_39;
  (* register *) pwire FA_cout_40;
  (* register *) pwire FA_cout_41;
  (* register *) pwire FA_cout_42;
  (* register *) pwire FA_cout_43;
  (* register *) pwire FA_cout_44;
  (* register *) pwire FA_cout_45;
  (* register *) pwire FA_cout_46;
  (* register *) pwire FA_cout_47;
  (* register *) pwire FA_cout_48;
  (* register *) pwire FA_cout_49;
  (* register *) pwire FA_cout_50;
  (* register *) pwire FA_cout_51;
  (* register *) pwire FA_cout_52;
  (* register *) pwire FA_cout_53;
  (* register *) pwire FA_cout_54;
  (* register *) pwire FA_cout_55;
  (* register *) pwire FA_cout_56;
  (* register *) pwire FA_cout_57;
  (* register *) pwire FA_cout_58;
  (* register *) pwire FA_cout_59;
  (* register *) pwire FA_cout_60;
  (* register *) pwire FA_cout_61;
  (* register *) pwire FA_cout_62;
  (* register *) pwire FA_cout_63;
  (* register *) pwire FA_cout_64;
  (* register *) pwire FA_cout_65;
  (* register *) pwire FA_cout_66;
  (* register *) pwire FA_cout_67;
  (* register *) pwire FA_cout_68;
  (* register *) pwire FA_cout_69;
  (* register *) pwire FA_cout_70;
  (* register *) pwire FA_cout_71;
  (* register *) pwire FA_cout_72;
  (* register *) pwire FA_cout_73;
  (* register *) pwire FA_cout_74;
  (* register *) pwire FA_cout_75;
  (* register *) pwire FA_cout_76;
  (* register *) pwire FA_cout_77;
  (* register *) pwire FA_cout_78;
  (* register *) pwire FA_cout_79;
  (* register *) pwire FA_cout_80;
  (* register *) pwire FA_cout_81;
  (* register *) pwire FA_cout_82;
  (* register *) pwire FA_cout_83;
  (* register *) pwire FA_cout_84;
  (* register *) pwire FA_cout_85;
  (* register *) pwire FA_cout_86;
  (* register *) pwire FA_cout_87;
  (* register *) pwire FA_cout_88;
  (* register *) pwire FA_cout_89;
  (* register *) pwire FA_cout_90;
  (* register *) pwire FA_cout_91;
  (* register *) pwire FA_cout_92;
  (* register *) pwire FA_cout_93;
  (* register *) pwire FA_cout_94;
  (* register *) pwire FA_cout_95;
  (* register *) pwire FA_cout_96;
  (* register *) pwire FA_cout_97;
  (* register *) pwire FA_cout_98;
  (* register *) pwire FA_cout_99;
  (* register *) pwire FA_cout_100;
  (* register *) pwire FA_cout_101;
  (* register *) pwire FA_cout_102;
  (* register *) pwire FA_cout_103;
  (* register *) pwire FA_cout_104;
  (* register *) pwire FA_cout_105;
  (* register *) pwire FA_cout_106;
  (* register *) pwire FA_cout_107;
  (* register *) pwire FA_cout_108;
  (* register *) pwire FA_cout_109;
  (* register *) pwire FA_cout_110;
  (* register *) pwire FA_cout_111;
  (* register *) pwire FA_cout_112;
  (* register *) pwire FA_cout_113;
  (* register *) pwire FA_cout_114;
  (* register *) pwire FA_cout_115;
  (* register *) pwire FA_cout_116;
  (* register *) pwire FA_cout_117;
  (* register *) pwire FA_cout_118;
  (* register *) pwire FA_cout_119;
  (* register *) pwire FA_cout_120;
  (* register *) pwire FA_cout_121;
  (* register *) pwire FA_cout_122;
  (* register *) pwire FA_cout_123;
  (* register *) pwire FA_cout_124;
  (* register *) pwire FA_cout_125;
  (* register *) pwire FA_cout_126;
  (* register *) pwire FA_cout_127;
  (* register *) pwire FA_cout_128;
  (* register *) pwire FA_cout_129;
  (* register *) pwire FA_cout_130;
  (* register *) pwire FA_cout_131;
  (* register *) pwire FA_cout_132;
  (* register *) pwire FA_cout_133;
  (* register *) pwire FA_cout_134;
  (* register *) pwire FA_cout_135;
  (* register *) pwire FA_cout_136;
  (* register *) pwire FA_cout_137;
  (* register *) pwire FA_cout_138;
  (* register *) pwire FA_cout_139;
  (* register *) pwire FA_cout_140;
  (* register *) pwire FA_cout_141;
  (* register *) pwire FA_cout_142;
  (* register *) pwire FA_cout_143;
  (* register *) pwire FA_cout_144;
  (* register *) pwire FA_cout_145;
  (* register *) pwire FA_cout_146;
  (* register *) pwire FA_cout_147;
  (* register *) pwire FA_cout_148;
  (* register *) pwire FA_cout_149;
  (* register *) pwire FA_cout_150;
  (* register *) pwire FA_cout_151;
  (* register *) pwire FA_cout_152;
  (* register *) pwire FA_cout_153;
  (* register *) pwire FA_cout_154;
  (* register *) pwire FA_cout_155;
  (* register *) pwire FA_cout_156;
  (* register *) pwire FA_cout_157;
  (* register *) pwire FA_cout_158;
  (* register *) pwire FA_cout_159;
  (* register *) pwire FA_cout_160;
  (* register *) pwire FA_cout_161;
  (* register *) pwire FA_cout_162;
  (* register *) pwire FA_cout_163;
  (* register *) pwire FA_cout_164;
  (* register *) pwire FA_cout_165;
  (* register *) pwire FA_cout_166;
  (* register *) pwire FA_cout_167;
  (* register *) pwire FA_cout_168;
  (* register *) pwire FA_cout_169;
  (* register *) pwire FA_cout_170;
  (* register *) pwire FA_cout_171;
  (* register *) pwire FA_cout_172;
  (* register *) pwire FA_cout_173;
  (* register *) pwire FA_cout_174;
  (* register *) pwire FA_cout_175;
  (* register *) pwire FA_cout_176;
  (* register *) pwire FA_cout_177;
  (* register *) pwire FA_cout_178;
  (* register *) pwire FA_cout_179;
  (* register *) pwire FA_cout_180;
  (* register *) pwire FA_cout_181;
  (* register *) pwire FA_cout_182;
  (* register *) pwire FA_cout_183;
  (* register *) pwire FA_cout_184;
  (* register *) pwire FA_cout_185;
  (* register *) pwire FA_cout_186;
  (* register *) pwire FA_cout_187;
  (* register *) pwire FA_cout_188;
  (* register *) pwire FA_cout_189;
  (* register *) pwire FA_cout_190;
  (* register *) pwire FA_cout_191;
  (* register *) pwire FA_cout_192;
  (* register *) pwire FA_cout_193;
  (* register *) pwire FA_cout_194;
  (* register *) pwire FA_cout_195;
  (* register *) pwire FA_cout_196;
  (* register *) pwire FA_cout_197;
  (* register *) pwire FA_cout_198;
  (* register *) pwire FA_cout_199;
  (* register *) pwire FA_cout_200;
  (* register *) pwire FA_cout_201;
  (* register *) pwire FA_cout_202;
  (* register *) pwire FA_cout_203;
  (* register *) pwire FA_cout_204;
  (* register *) pwire FA_cout_205;
  (* register *) pwire FA_cout_206;
  (* register *) pwire FA_cout_207;
  (* register *) pwire FA_cout_208;
  (* register *) pwire FA_cout_209;
  (* register *) pwire FA_cout_210;
  (* register *) pwire FA_cout_211;
  (* register *) pwire FA_cout_212;
  (* register *) pwire FA_cout_213;
  (* register *) pwire FA_cout_214;
  (* register *) pwire FA_cout_215;
  (* register *) pwire FA_cout_216;
  (* register *) pwire FA_cout_217;
  (* register *) pwire FA_cout_218;
  (* register *) pwire FA_cout_219;
  (* register *) pwire FA_cout_220;
  (* register *) pwire FA_cout_221;
  (* register *) pwire FA_cout_222;
  (* register *) pwire FA_cout_223;
  (* register *) pwire FA_cout_224;
  (* register *) pwire FA_cout_225;
  (* register *) pwire FA_cout_226;
  (* register *) pwire FA_cout_227;
  (* register *) pwire FA_cout_228;
  (* register *) pwire FA_cout_229;
  (* register *) pwire FA_cout_230;
  (* register *) pwire FA_cout_231;
  (* register *) pwire FA_cout_232;
  (* register *) pwire FA_cout_233;
  (* register *) pwire FA_cout_234;
  (* register *) pwire FA_cout_235;
  (* register *) pwire FA_cout_236;
  (* register *) pwire FA_cout_237;
  (* register *) pwire FA_cout_238;
  (* register *) pwire FA_cout_239;
  (* register *) pwire FA_cout_240;
  (* register *) pwire FA_cout_241;
  (* register *) pwire FA_cout_242;
  (* register *) pwire FA_cout_243;
  (* register *) pwire FA_cout_244;
  (* register *) pwire FA_cout_245;
  (* register *) pwire FA_cout_246;
  (* register *) pwire FA_cout_247;
  (* register *) pwire FA_cout_248;
  (* register *) pwire FA_cout_249;
  (* register *) pwire FA_cout_250;
  (* register *) pwire FA_cout_251;
  (* register *) pwire FA_cout_252;
  (* register *) pwire FA_cout_253;
  (* register *) pwire FA_cout_254;
  (* register *) pwire FA_cout_255;
  (* register *) pwire FA_cout_256;
  (* register *) pwire FA_cout_257;
  (* register *) pwire FA_cout_258;
  (* register *) pwire FA_cout_259;
  (* register *) pwire FA_cout_260;
  (* register *) pwire FA_cout_261;
  (* register *) pwire FA_cout_262;
  (* register *) pwire FA_cout_263;
  (* register *) pwire FA_cout_264;
  (* register *) pwire FA_cout_265;
  (* register *) pwire FA_cout_266;
  (* register *) pwire FA_cout_267;
  (* register *) pwire FA_cout_268;
  (* register *) pwire FA_cout_269;
  (* register *) pwire FA_cout_270;
  (* register *) pwire FA_cout_271;
  (* register *) pwire FA_cout_272;
  (* register *) pwire FA_cout_273;
  (* register *) pwire FA_cout_274;
  (* register *) pwire FA_cout_275;
  (* register *) pwire FA_cout_276;
  (* register *) pwire FA_cout_277;
  (* register *) pwire FA_cout_278;
  (* register *) pwire FA_cout_279;
  (* register *) pwire FA_cout_280;
  (* register *) pwire FA_cout_281;
  (* register *) pwire FA_cout_282;
  (* register *) pwire FA_cout_283;
  (* register *) pwire FA_cout_284;
  (* register *) pwire FA_cout_285;
  (* register *) pwire FA_cout_286;
  (* register *) pwire FA_cout_287;
  (* register *) pwire FA_cout_288;
  (* register *) pwire FA_cout_289;
  (* register *) pwire FA_cout_290;
  (* register *) pwire FA_cout_291;
  (* register *) pwire FA_cout_292;
  (* register *) pwire FA_cout_293;
  (* register *) pwire FA_cout_294;
  (* register *) pwire FA_cout_295;
  (* register *) pwire FA_cout_296;
  (* register *) pwire FA_cout_297;
  (* register *) pwire FA_cout_298;
  (* register *) pwire FA_cout_299;
  (* register *) pwire FA_cout_300;
  (* register *) pwire FA_cout_301;
  (* register *) pwire FA_cout_302;
  (* register *) pwire FA_cout_303;
  (* register *) pwire FA_cout_304;
  (* register *) pwire FA_cout_305;
  (* register *) pwire FA_cout_306;
  (* register *) pwire FA_cout_307;
  (* register *) pwire FA_cout_308;
  (* register *) pwire FA_cout_309;
  (* register *) pwire FA_cout_310;
  (* register *) pwire FA_cout_311;
  (* register *) pwire FA_cout_312;
  (* register *) pwire FA_cout_313;
  (* register *) pwire FA_cout_314;
  (* register *) pwire FA_cout_315;
  (* register *) pwire FA_cout_316;
  (* register *) pwire FA_cout_317;
  (* register *) pwire FA_cout_318;
  (* register *) pwire FA_cout_319;
  (* register *) pwire FA_cout_320;
  (* register *) pwire FA_cout_321;
  (* register *) pwire FA_cout_322;
  (* register *) pwire FA_cout_323;
  (* register *) pwire FA_cout_324;
  (* register *) pwire FA_cout_325;
  (* register *) pwire FA_cout_326;
  (* register *) pwire FA_cout_327;
  (* register *) pwire FA_cout_328;
  (* register *) pwire FA_cout_329;
  (* register *) pwire FA_cout_330;
  (* register *) pwire FA_cout_331;
  (* register *) pwire FA_cout_332;
  (* register *) pwire FA_cout_333;
  (* register *) pwire FA_cout_334;
  (* register *) pwire FA_cout_335;
  (* register *) pwire FA_cout_336;
  (* register *) pwire FA_cout_337;
  (* register *) pwire FA_cout_338;
  (* register *) pwire FA_cout_339;
  (* register *) pwire FA_cout_340;
  (* register *) pwire FA_cout_341;
  (* register *) pwire FA_cout_342;
  (* register *) pwire FA_cout_343;
  (* register *) pwire FA_cout_344;
  (* register *) pwire FA_cout_345;
  (* register *) pwire FA_cout_346;
  (* register *) pwire FA_cout_347;
  (* register *) pwire FA_cout_348;
  (* register *) pwire FA_cout_349;
  (* register *) pwire FA_cout_350;
  (* register *) pwire FA_cout_351;
  (* register *) pwire FA_cout_352;
  (* register *) pwire FA_cout_353;
  (* register *) pwire FA_cout_354;
  (* register *) pwire FA_cout_355;
  (* register *) pwire FA_cout_356;
  (* register *) pwire FA_cout_357;
  (* register *) pwire FA_cout_358;
  (* register *) pwire FA_cout_359;
  (* register *) pwire FA_cout_360;
  (* register *) pwire FA_cout_361;
  (* register *) pwire FA_cout_362;
  (* register *) pwire FA_cout_363;
  (* register *) pwire FA_cout_364;
  (* register *) pwire FA_cout_365;
  (* register *) pwire FA_cout_366;
  (* register *) pwire FA_cout_367;
  (* register *) pwire FA_cout_368;
  (* register *) pwire FA_cout_369;
  (* register *) pwire FA_cout_370;
  (* register *) pwire FA_cout_371;
  (* register *) pwire FA_cout_372;
  (* register *) pwire FA_cout_373;
  (* register *) pwire FA_cout_374;
  (* register *) pwire FA_cout_375;
  (* register *) pwire FA_cout_376;
  (* register *) pwire FA_cout_377;
  (* register *) pwire FA_cout_378;
  (* register *) pwire FA_cout_379;
  (* register *) pwire FA_cout_380;
  (* register *) pwire FA_cout_381;
  (* register *) pwire FA_cout_382;
  (* register *) pwire FA_cout_383;
  (* register *) pwire FA_cout_384;
  (* register *) pwire FA_cout_385;
  (* register *) pwire FA_cout_386;
  (* register *) pwire FA_cout_387;
  (* register *) pwire FA_cout_388;
  (* register *) pwire FA_cout_389;
  (* register *) pwire FA_cout_390;
  (* register *) pwire FA_cout_391;
  (* register *) pwire FA_cout_392;
  (* register *) pwire FA_cout_393;
  (* register *) pwire FA_cout_394;
  (* register *) pwire FA_cout_395;
  (* register *) pwire FA_cout_396;
  (* register *) pwire FA_cout_397;
  (* register *) pwire FA_cout_398;
  (* register *) pwire FA_cout_399;
  (* register *) pwire FA_cout_400;
  (* register *) pwire FA_cout_401;
  (* register *) pwire FA_cout_402;
  (* register *) pwire FA_cout_403;
  (* register *) pwire FA_cout_404;
  (* register *) pwire FA_cout_405;
  (* register *) pwire FA_cout_406;
  (* register *) pwire FA_cout_407;
  (* register *) pwire FA_cout_408;
  (* register *) pwire FA_cout_409;
  (* register *) pwire FA_cout_410;
  (* register *) pwire FA_cout_411;
  (* register *) pwire FA_cout_412;
  (* register *) pwire FA_cout_413;
  (* register *) pwire FA_cout_414;
  (* register *) pwire FA_cout_415;
  (* register *) pwire FA_cout_416;
  (* register *) pwire FA_cout_417;
  (* register *) pwire FA_cout_418;
  (* register *) pwire FA_cout_419;
  (* register *) pwire FA_cout_420;
  (* register *) pwire FA_cout_421;
  (* register *) pwire FA_cout_422;
  (* register *) pwire FA_cout_423;
  (* register *) pwire FA_cout_424;
  (* register *) pwire FA_cout_425;
  (* register *) pwire FA_cout_426;
  (* register *) pwire FA_cout_427;
  (* register *) pwire FA_cout_428;
  (* register *) pwire FA_cout_429;
  (* register *) pwire FA_cout_430;
  (* register *) pwire FA_cout_431;
  (* register *) pwire FA_cout_432;
  (* register *) pwire FA_cout_433;
  (* register *) pwire FA_cout_434;
  (* register *) pwire FA_cout_435;
  (* register *) pwire FA_cout_436;
  (* register *) pwire FA_cout_437;
  (* register *) pwire FA_cout_438;
  (* register *) pwire FA_cout_439;
  (* register *) pwire FA_cout_440;
  (* register *) pwire FA_cout_441;
  (* register *) pwire FA_cout_442;
  (* register *) pwire FA_cout_443;
  (* register *) pwire FA_cout_444;
  (* register *) pwire FA_cout_445;
  (* register *) pwire FA_cout_446;
  (* register *) pwire FA_cout_447;
  (* register *) pwire FA_cout_448;
  (* register *) pwire FA_cout_449;
  (* register *) pwire FA_cout_450;
  (* register *) pwire FA_cout_451;
  (* register *) pwire FA_cout_452;
  (* register *) pwire FA_cout_453;
  (* register *) pwire FA_cout_454;
  (* register *) pwire FA_cout_455;
  (* register *) pwire FA_cout_456;
  (* register *) pwire FA_cout_457;
  (* register *) pwire FA_cout_458;
  (* register *) pwire FA_cout_459;
  (* register *) pwire FA_cout_460;
  (* register *) pwire FA_cout_461;
  (* register *) pwire FA_cout_462;
  (* register *) pwire FA_cout_463;
  (* register *) pwire FA_cout_464;
  (* register *) pwire FA_cout_465;
  (* register *) pwire FA_cout_466;
  (* register *) pwire FA_cout_467;
  (* register *) pwire FA_cout_468;
  (* register *) pwire FA_cout_469;
  (* register *) pwire FA_cout_470;
  (* register *) pwire FA_cout_471;
  (* register *) pwire FA_cout_472;
  (* register *) pwire FA_cout_473;
  (* register *) pwire FA_cout_474;
  (* register *) pwire FA_cout_475;
  (* register *) pwire FA_cout_476;
  (* register *) pwire FA_cout_477;
  (* register *) pwire FA_cout_478;
  (* register *) pwire FA_cout_479;
  (* register *) pwire FA_cout_480;
  (* register *) pwire FA_cout_481;
  (* register *) pwire FA_cout_482;
  (* register *) pwire FA_cout_483;
  (* register *) pwire HA_out_0;
  (* register *) pwire HA_out_1;
  (* register *) pwire HA_out_2;
  (* register *) pwire HA_out_3;
  (* register *) pwire HA_out_4;
  (* register *) pwire HA_out_5;
  (* register *) pwire HA_out_6;
  (* register *) pwire HA_out_7;
  (* register *) pwire HA_out_8;
  (* register *) pwire HA_out_9;
  (* register *) pwire HA_out_10;
  (* register *) pwire HA_out_11;
  (* register *) pwire HA_out_12;
  (* register *) pwire HA_out_13;
  (* register *) pwire HA_out_14;
  (* register *) pwire HA_out_15;
  (* register *) pwire HA_out_16;
  (* register *) pwire HA_out_17;
  (* register *) pwire HA_out_18;
  (* register *) pwire HA_out_19;
  (* register *) pwire HA_out_20;
  (* register *) pwire HA_out_21;
  (* register *) pwire HA_out_22;
  (* register *) pwire HA_out_23;
  (* register *) pwire HA_out_24;
  (* register *) pwire HA_out_25;
  (* register *) pwire HA_out_26;
  (* register *) pwire HA_out_27;
  (* register *) pwire HA_out_28;
  (* register *) pwire HA_out_29;
  (* register *) pwire HA_out_30;
  (* register *) pwire HA_out_31;
  (* register *) pwire HA_out_32;
  (* register *) pwire HA_out_33;
  (* register *) pwire HA_out_34;
  (* register *) pwire HA_out_35;
  (* register *) pwire HA_out_36;
  (* register *) pwire HA_out_37;
  (* register *) pwire HA_out_38;
  (* register *) pwire HA_out_39;
  (* register *) pwire HA_out_40;
  (* register *) pwire HA_out_41;
  (* register *) pwire HA_out_42;
  (* register *) pwire HA_out_43;
  (* register *) pwire HA_out_44;
  (* register *) pwire HA_out_45;
  (* register *) pwire HA_out_46;
  (* register *) pwire HA_out_47;
  (* register *) pwire HA_out_48;
  (* register *) pwire HA_out_49;
  (* register *) pwire HA_out_50;
  (* register *) pwire HA_out_51;
  (* register *) pwire HA_out_52;
  (* register *) pwire HA_out_53;
  (* register *) pwire HA_out_54;
  (* register *) pwire HA_out_55;
  (* register *) pwire HA_out_56;
  (* register *) pwire HA_out_57;
  (* register *) pwire HA_out_58;
  (* register *) pwire HA_out_59;
  (* register *) pwire HA_out_60;
  (* register *) pwire HA_out_61;
  (* register *) pwire HA_out_62;
  (* register *) pwire HA_out_63;
  (* register *) pwire HA_out_64;
  (* register *) pwire HA_out_65;
  (* register *) pwire HA_out_66;
  (* register *) pwire HA_out_67;
  (* register *) pwire HA_out_68;
  (* register *) pwire HA_out_69;
  (* register *) pwire HA_out_70;
  (* register *) pwire HA_out_71;
  (* register *) pwire HA_out_72;
  (* register *) pwire HA_out_73;
  (* register *) pwire HA_out_74;
  (* register *) pwire HA_out_75;
  (* register *) pwire HA_out_76;
  (* register *) pwire HA_out_77;
  (* register *) pwire HA_out_78;
  (* register *) pwire HA_out_79;
  (* register *) pwire HA_out_80;
  (* register *) pwire HA_out_81;
  (* register *) pwire HA_out_82;
  (* register *) pwire HA_out_83;
  (* register *) pwire HA_out_84;
  (* register *) pwire HA_out_85;
  (* register *) pwire HA_out_86;
  (* register *) pwire HA_out_87;
  (* register *) pwire HA_out_88;
  (* register *) pwire HA_out_89;
  (* register *) pwire HA_out_90;
  (* register *) pwire HA_out_91;
  (* register *) pwire HA_out_92;
  (* register *) pwire HA_out_93;
  (* register *) pwire HA_out_94;
  (* register *) pwire HA_out_95;
  (* register *) pwire HA_out_96;
  (* register *) pwire HA_out_97;
  (* register *) pwire HA_out_98;
  (* register *) pwire HA_out_99;
  (* register *) pwire HA_out_100;
  (* register *) pwire HA_out_101;
  (* register *) pwire HA_out_102;
  (* register *) pwire HA_out_103;
  (* register *) pwire HA_out_104;
  (* register *) pwire HA_out_105;
  (* register *) pwire HA_out_106;
  (* register *) pwire HA_out_107;
  (* register *) pwire HA_out_108;
  (* register *) pwire HA_out_109;
  (* register *) pwire HA_out_110;
  (* register *) pwire HA_out_111;
  (* register *) pwire HA_out_112;
  (* register *) pwire HA_out_113;
  (* register *) pwire HA_out_114;
  (* register *) pwire HA_out_115;
  (* register *) pwire HA_out_116;
  (* register *) pwire HA_out_117;
  (* register *) pwire HA_out_118;
  (* register *) pwire HA_out_119;
  (* register *) pwire HA_out_120;
  (* register *) pwire HA_out_121;
  (* register *) pwire HA_out_122;
  (* register *) pwire HA_out_123;
  (* register *) pwire HA_out_124;
  (* register *) pwire HA_out_125;
  (* register *) pwire HA_out_126;
  (* register *) pwire HA_out_127;
  (* register *) pwire HA_out_128;
  (* register *) pwire HA_out_129;
  (* register *) pwire HA_out_130;
  (* register *) pwire HA_out_131;
  (* register *) pwire HA_out_132;
  (* register *) pwire HA_out_133;
  (* register *) pwire HA_out_134;
  (* register *) pwire HA_out_135;
  (* register *) pwire HA_out_136;
  (* register *) pwire HA_out_137;
  (* register *) pwire HA_out_138;
  (* register *) pwire HA_cout_0;
  (* register *) pwire HA_cout_1;
  (* register *) pwire HA_cout_2;
  (* register *) pwire HA_cout_3;
  (* register *) pwire HA_cout_4;
  (* register *) pwire HA_cout_5;
  (* register *) pwire HA_cout_6;
  (* register *) pwire HA_cout_7;
  (* register *) pwire HA_cout_8;
  (* register *) pwire HA_cout_9;
  (* register *) pwire HA_cout_10;
  (* register *) pwire HA_cout_11;
  (* register *) pwire HA_cout_12;
  (* register *) pwire HA_cout_13;
  (* register *) pwire HA_cout_14;
  (* register *) pwire HA_cout_15;
  (* register *) pwire HA_cout_16;
  (* register *) pwire HA_cout_17;
  (* register *) pwire HA_cout_18;
  (* register *) pwire HA_cout_19;
  (* register *) pwire HA_cout_20;
  (* register *) pwire HA_cout_21;
  (* register *) pwire HA_cout_22;
  (* register *) pwire HA_cout_23;
  (* register *) pwire HA_cout_24;
  (* register *) pwire HA_cout_25;
  (* register *) pwire HA_cout_26;
  (* register *) pwire HA_cout_27;
  (* register *) pwire HA_cout_28;
  (* register *) pwire HA_cout_29;
  (* register *) pwire HA_cout_30;
  (* register *) pwire HA_cout_31;
  (* register *) pwire HA_cout_32;
  (* register *) pwire HA_cout_33;
  (* register *) pwire HA_cout_34;
  (* register *) pwire HA_cout_35;
  (* register *) pwire HA_cout_36;
  (* register *) pwire HA_cout_37;
  (* register *) pwire HA_cout_38;
  (* register *) pwire HA_cout_39;
  (* register *) pwire HA_cout_40;
  (* register *) pwire HA_cout_41;
  (* register *) pwire HA_cout_42;
  (* register *) pwire HA_cout_43;
  (* register *) pwire HA_cout_44;
  (* register *) pwire HA_cout_45;
  (* register *) pwire HA_cout_46;
  (* register *) pwire HA_cout_47;
  (* register *) pwire HA_cout_48;
  (* register *) pwire HA_cout_49;
  (* register *) pwire HA_cout_50;
  (* register *) pwire HA_cout_51;
  (* register *) pwire HA_cout_52;
  (* register *) pwire HA_cout_53;
  (* register *) pwire HA_cout_54;
  (* register *) pwire HA_cout_55;
  (* register *) pwire HA_cout_56;
  (* register *) pwire HA_cout_57;
  (* register *) pwire HA_cout_58;
  (* register *) pwire HA_cout_59;
  (* register *) pwire HA_cout_60;
  (* register *) pwire HA_cout_61;
  (* register *) pwire HA_cout_62;
  (* register *) pwire HA_cout_63;
  (* register *) pwire HA_cout_64;
  (* register *) pwire HA_cout_65;
  (* register *) pwire HA_cout_66;
  (* register *) pwire HA_cout_67;
  (* register *) pwire HA_cout_68;
  (* register *) pwire HA_cout_69;
  (* register *) pwire HA_cout_70;
  (* register *) pwire HA_cout_71;
  (* register *) pwire HA_cout_72;
  (* register *) pwire HA_cout_73;
  (* register *) pwire HA_cout_74;
  (* register *) pwire HA_cout_75;
  (* register *) pwire HA_cout_76;
  (* register *) pwire HA_cout_77;
  (* register *) pwire HA_cout_78;
  (* register *) pwire HA_cout_79;
  (* register *) pwire HA_cout_80;
  (* register *) pwire HA_cout_81;
  (* register *) pwire HA_cout_82;
  (* register *) pwire HA_cout_83;
  (* register *) pwire HA_cout_84;
  (* register *) pwire HA_cout_85;
  (* register *) pwire HA_cout_86;
  (* register *) pwire HA_cout_87;
  (* register *) pwire HA_cout_88;
  (* register *) pwire HA_cout_89;
  (* register *) pwire HA_cout_90;
  (* register *) pwire HA_cout_91;
  (* register *) pwire HA_cout_92;
  (* register *) pwire HA_cout_93;
  (* register *) pwire HA_cout_94;
  (* register *) pwire HA_cout_95;
  (* register *) pwire HA_cout_96;
  (* register *) pwire HA_cout_97;
  (* register *) pwire HA_cout_98;
  (* register *) pwire HA_cout_99;
  (* register *) pwire HA_cout_100;
  (* register *) pwire HA_cout_101;
  (* register *) pwire HA_cout_102;
  (* register *) pwire HA_cout_103;
  (* register *) pwire HA_cout_104;
  (* register *) pwire HA_cout_105;
  (* register *) pwire HA_cout_106;
  (* register *) pwire HA_cout_107;
  (* register *) pwire HA_cout_108;
  (* register *) pwire HA_cout_109;
  (* register *) pwire HA_cout_110;
  (* register *) pwire HA_cout_111;
  (* register *) pwire HA_cout_112;
  (* register *) pwire HA_cout_113;
  (* register *) pwire HA_cout_114;
  (* register *) pwire HA_cout_115;
  (* register *) pwire HA_cout_116;
  (* register *) pwire HA_cout_117;
  (* register *) pwire HA_cout_118;
  (* register *) pwire HA_cout_119;
  (* register *) pwire HA_cout_120;
  (* register *) pwire HA_cout_121;
  (* register *) pwire HA_cout_122;
  (* register *) pwire HA_cout_123;
  (* register *) pwire HA_cout_124;
  (* register *) pwire HA_cout_125;
  (* register *) pwire HA_cout_126;
  (* register *) pwire HA_cout_127;
  (* register *) pwire HA_cout_128;
  (* register *) pwire HA_cout_129;
  (* register *) pwire HA_cout_130;
  (* register *) pwire HA_cout_131;
  (* register *) pwire HA_cout_132;
  (* register *) pwire HA_cout_133;
  (* register *) pwire HA_cout_134;
  (* register *) pwire HA_cout_135;
  (* register *) pwire HA_cout_136;
  (* register *) pwire HA_cout_137;
  (* register *) pwire HA_cout_138;
  (* register *) pwire [23:0] inp_0;

  (* register *) pwire [23:0] inp_1;

  (* register *) pwire [23:0] inp_2;

  (* register *) pwire [23:0] inp_3;

  (* register *) pwire [23:0] inp_4;

  (* register *) pwire [23:0] inp_5;

  (* register *) pwire [23:0] inp_6;

  (* register *) pwire [23:0] inp_7;

  (* register *) pwire [23:0] inp_8;

  (* register *) pwire [23:0] inp_9;

  (* register *) pwire [23:0] inp_10;

  (* register *) pwire [23:0] inp_11;

  (* register *) pwire [23:0] inp_12;

  (* register *) pwire [23:0] inp_13;

  (* register *) pwire [23:0] inp_14;

  (* register *) pwire [23:0] inp_15;

  (* register *) pwire [23:0] inp_16;

  (* register *) pwire [23:0] inp_17;

  (* register *) pwire [23:0] inp_18;

  (* register *) pwire [23:0] inp_19;

  (* register *) pwire [23:0] inp_20;

  (* register *) pwire [23:0] inp_21;

  (* register *) pwire [23:0] inp_22;

  (* register *) pwire [23:0] inp_23;

  assign inp_0=C & {24{R[0]}};
  assign inp_1=C & {24{R[1]}};
  assign inp_2=C & {24{R[2]}};
  assign inp_3=C & {24{R[3]}};
  assign inp_4=C & {24{R[4]}};
  assign inp_5=C & {24{R[5]}};
  assign inp_6=C & {24{R[6]}};
  assign inp_7=C & {24{R[7]}};
  assign inp_8=C & {24{R[8]}};
  assign inp_9=C & {24{R[9]}};
  assign inp_10=C & {24{R[10]}};
  assign inp_11=C & {24{R[11]}};
  assign inp_12=C & {24{R[12]}};
  assign inp_13=C & {24{R[13]}};
  assign inp_14=C & {24{R[14]}};
  assign inp_15=C & {24{R[15]}};
  assign inp_16=C & {24{R[16]}};
  assign inp_17=C & {24{R[17]}};
  assign inp_18=C & {24{R[18]}};
  assign inp_19=C & {24{R[19]}};
  assign inp_20=C & {24{R[20]}};
  assign inp_21=C & {24{R[21]}};
  assign inp_22=C & {24{R[22]}};
  assign inp_23=C & {24{R[23]}};
  assign A_out[0]=REGS_283;
  assign A_out[1]=REGS_284;
  assign A_out[2]=REGS_285;
  assign A_out[3]=REGS_286;
  assign A_out[4]=REGS_287;
  assign A_out[5]=REGS_288;
  assign A_out[6]=REGS_289;
  assign A_out[7]=HA_out_105;
  assign A_out[8]=HA_cout_105;
  assign A_out[9]=HA_cout_106;
  assign A_out[10]=HA_cout_107;
  assign A_out[11]=HA_cout_108;
  assign A_out[12]=HA_cout_109;
  assign A_out[13]=HA_cout_110;
  assign A_out[14]=HA_cout_111;
  assign A_out[15]=HA_cout_112;
  assign A_out[16]=HA_cout_113;
  assign A_out[17]=HA_cout_114;
  assign A_out[18]=HA_cout_115;
  assign A_out[19]=HA_cout_116;
  assign A_out[20]=HA_cout_117;
  assign A_out[21]=HA_cout_118;
  assign A_out[22]=HA_cout_119;
  assign A_out[23]=FA_cout_476;
  assign A_out[24]=FA_cout_477;
  assign A_out[25]=FA_cout_478;
  assign A_out[26]=FA_cout_479;
  assign A_out[27]=FA_cout_480;
  assign A_out[28]=FA_cout_481;
  assign A_out[29]=FA_cout_482;
  assign A_out[30]=FA_cout_483;
  assign B_out[8]=HA_out_106;
  assign B_out[9]=HA_out_107;
  assign B_out[10]=HA_out_108;
  assign B_out[11]=HA_out_109;
  assign B_out[12]=HA_out_110;
  assign B_out[13]=HA_out_111;
  assign B_out[14]=HA_out_112;
  assign B_out[15]=HA_out_113;
  assign B_out[16]=HA_out_114;
  assign B_out[17]=HA_out_115;
  assign B_out[18]=HA_out_116;
  assign B_out[19]=HA_out_117;
  assign B_out[20]=HA_out_118;
  assign B_out[21]=HA_out_119;
  assign B_out[22]=FA_out_476;
  assign B_out[23]=FA_out_477;
  assign B_out[24]=FA_out_478;
  assign B_out[25]=FA_out_479;
  assign B_out[26]=FA_out_480;
  assign B_out[27]=FA_out_481;
  assign B_out[28]=FA_out_482;
  assign B_out[29]=FA_out_483;
  assign B_out[30]=HA_out_120;
  assign A_out[31]=HA_cout_120;
  assign B_out[31]=HA_out_121;
  assign A_out[32]=HA_cout_121;
  assign B_out[32]=HA_out_122;
  assign A_out[33]=HA_cout_122;
  assign B_out[33]=HA_out_123;
  assign A_out[34]=HA_cout_123;
  assign B_out[34]=HA_out_124;
  assign A_out[35]=HA_cout_124;
  assign B_out[35]=HA_out_125;
  assign A_out[36]=HA_cout_125;
  assign B_out[36]=HA_out_126;
  assign A_out[37]=HA_cout_126;
  assign B_out[37]=HA_out_127;
  assign A_out[38]=HA_cout_127;
  assign B_out[38]=HA_out_128;
  assign A_out[39]=HA_cout_128;
  assign B_out[39]=HA_out_129;
  assign A_out[40]=HA_cout_129;
  assign B_out[40]=HA_out_130;
  assign A_out[41]=HA_cout_130;
  assign B_out[41]=HA_out_131;
  assign A_out[42]=HA_cout_131;
  assign B_out[42]=HA_out_132;
  assign A_out[43]=HA_cout_132;
  assign B_out[43]=HA_out_133;
  assign A_out[44]=HA_cout_133;
  assign B_out[44]=HA_out_134;
  assign A_out[45]=HA_cout_134;
  assign B_out[45]=HA_out_135;
  assign A_out[46]=HA_cout_135;
  assign B_out[46]=HA_out_136;
  assign A_out[47]=HA_cout_136;
  assign B_out[47]=HA_out_137;
  assign B_out[0]=1'b0;
  assign B_out[1]=1'b0;
  assign B_out[2]=1'b0;
  assign B_out[3]=1'b0;
  assign B_out[4]=1'b0;
  assign B_out[5]=1'b0;
  assign B_out[6]=1'b0;
  assign B_out[7]=1'b0;

  assign {FA_cout_0,FA_out_0}=inp_0[2]+inp_1[1]+inp_2[0];
  assign {FA_cout_1,FA_out_1}=inp_0[3]+inp_1[2]+inp_2[1];
  assign {FA_cout_2,FA_out_2}=inp_0[4]+inp_1[3]+inp_2[2];
  assign {FA_cout_3,FA_out_3}=inp_0[5]+inp_1[4]+inp_2[3];
  assign {FA_cout_4,FA_out_4}=inp_0[6]+inp_1[5]+inp_2[4];
  assign {FA_cout_5,FA_out_5}=inp_0[7]+inp_1[6]+inp_2[5];
  assign {FA_cout_6,FA_out_6}=inp_0[8]+inp_1[7]+inp_2[6];
  assign {FA_cout_7,FA_out_7}=inp_0[9]+inp_1[8]+inp_2[7];
  assign {FA_cout_8,FA_out_8}=inp_0[10]+inp_1[9]+inp_2[8];
  assign {FA_cout_9,FA_out_9}=inp_0[11]+inp_1[10]+inp_2[9];
  assign {FA_cout_10,FA_out_10}=inp_0[12]+inp_1[11]+inp_2[10];
  assign {FA_cout_11,FA_out_11}=inp_0[13]+inp_1[12]+inp_2[11];
  assign {FA_cout_12,FA_out_12}=inp_0[14]+inp_1[13]+inp_2[12];
  assign {FA_cout_13,FA_out_13}=inp_0[15]+inp_1[14]+inp_2[13];
  assign {FA_cout_14,FA_out_14}=inp_0[16]+inp_1[15]+inp_2[14];
  assign {FA_cout_15,FA_out_15}=inp_0[17]+inp_1[16]+inp_2[15];
  assign {FA_cout_16,FA_out_16}=inp_0[18]+inp_1[17]+inp_2[16];
  assign {FA_cout_17,FA_out_17}=inp_0[19]+inp_1[18]+inp_2[17];
  assign {FA_cout_18,FA_out_18}=inp_0[20]+inp_1[19]+inp_2[18];
  assign {FA_cout_19,FA_out_19}=inp_0[21]+inp_1[20]+inp_2[19];
  assign {FA_cout_20,FA_out_20}=inp_0[22]+inp_1[21]+inp_2[20];
  assign {FA_cout_21,FA_out_21}=inp_0[23]+inp_1[22]+inp_2[21];
  assign {FA_cout_22,FA_out_22}=inp_1[23]+inp_2[22]+inp_3[21];
  assign {FA_cout_23,FA_out_23}=inp_2[23]+inp_3[22]+inp_4[21];
  assign {FA_cout_24,FA_out_24}=inp_3[2]+inp_4[1]+inp_5[0];
  assign {FA_cout_25,FA_out_25}=inp_3[3]+inp_4[2]+inp_5[1];
  assign {FA_cout_26,FA_out_26}=inp_3[4]+inp_4[3]+inp_5[2];
  assign {FA_cout_27,FA_out_27}=inp_3[5]+inp_4[4]+inp_5[3];
  assign {FA_cout_28,FA_out_28}=inp_3[6]+inp_4[5]+inp_5[4];
  assign {FA_cout_29,FA_out_29}=inp_3[7]+inp_4[6]+inp_5[5];
  assign {FA_cout_30,FA_out_30}=inp_3[8]+inp_4[7]+inp_5[6];
  assign {FA_cout_31,FA_out_31}=inp_3[9]+inp_4[8]+inp_5[7];
  assign {FA_cout_32,FA_out_32}=inp_3[10]+inp_4[9]+inp_5[8];
  assign {FA_cout_33,FA_out_33}=inp_3[11]+inp_4[10]+inp_5[9];
  assign {FA_cout_34,FA_out_34}=inp_3[12]+inp_4[11]+inp_5[10];
  assign {FA_cout_35,FA_out_35}=inp_3[13]+inp_4[12]+inp_5[11];
  assign {FA_cout_36,FA_out_36}=inp_3[14]+inp_4[13]+inp_5[12];
  assign {FA_cout_37,FA_out_37}=inp_3[15]+inp_4[14]+inp_5[13];
  assign {FA_cout_38,FA_out_38}=inp_3[16]+inp_4[15]+inp_5[14];
  assign {FA_cout_39,FA_out_39}=inp_3[17]+inp_4[16]+inp_5[15];
  assign {FA_cout_40,FA_out_40}=inp_3[18]+inp_4[17]+inp_5[16];
  assign {FA_cout_41,FA_out_41}=inp_3[19]+inp_4[18]+inp_5[17];
  assign {FA_cout_42,FA_out_42}=inp_3[20]+inp_4[19]+inp_5[18];
  assign {FA_cout_43,FA_out_43}=inp_3[23]+inp_4[22]+inp_5[21];
  assign {FA_cout_44,FA_out_44}=inp_4[20]+inp_5[19]+inp_6[18];
  assign {FA_cout_45,FA_out_45}=inp_4[23]+inp_5[22]+inp_6[21];
  assign {FA_cout_46,FA_out_46}=inp_5[20]+inp_6[19]+inp_7[18];
  assign {FA_cout_47,FA_out_47}=inp_5[23]+inp_6[22]+inp_7[21];
  assign {FA_cout_48,FA_out_48}=inp_6[2]+inp_7[1]+inp_8[0];
  assign {FA_cout_49,FA_out_49}=inp_6[3]+inp_7[2]+inp_8[1];
  assign {FA_cout_50,FA_out_50}=inp_6[4]+inp_7[3]+inp_8[2];
  assign {FA_cout_51,FA_out_51}=inp_6[5]+inp_7[4]+inp_8[3];
  assign {FA_cout_52,FA_out_52}=inp_6[6]+inp_7[5]+inp_8[4];
  assign {FA_cout_53,FA_out_53}=inp_6[7]+inp_7[6]+inp_8[5];
  assign {FA_cout_54,FA_out_54}=inp_6[8]+inp_7[7]+inp_8[6];
  assign {FA_cout_55,FA_out_55}=inp_6[9]+inp_7[8]+inp_8[7];
  assign {FA_cout_56,FA_out_56}=inp_6[10]+inp_7[9]+inp_8[8];
  assign {FA_cout_57,FA_out_57}=inp_6[11]+inp_7[10]+inp_8[9];
  assign {FA_cout_58,FA_out_58}=inp_6[12]+inp_7[11]+inp_8[10];
  assign {FA_cout_59,FA_out_59}=inp_6[13]+inp_7[12]+inp_8[11];
  assign {FA_cout_60,FA_out_60}=inp_6[14]+inp_7[13]+inp_8[12];
  assign {FA_cout_61,FA_out_61}=inp_6[15]+inp_7[14]+inp_8[13];
  assign {FA_cout_62,FA_out_62}=inp_6[16]+inp_7[15]+inp_8[14];
  assign {FA_cout_63,FA_out_63}=inp_6[17]+inp_7[16]+inp_8[15];
  assign {FA_cout_64,FA_out_64}=inp_6[20]+inp_7[19]+inp_8[18];
  assign {FA_cout_65,FA_out_65}=inp_6[23]+inp_7[22]+inp_8[21];
  assign {FA_cout_66,FA_out_66}=inp_7[17]+inp_8[16]+inp_9[15];
  assign {FA_cout_67,FA_out_67}=inp_7[20]+inp_8[19]+inp_9[18];
  assign {FA_cout_68,FA_out_68}=inp_7[23]+inp_8[22]+inp_9[21];
  assign {FA_cout_69,FA_out_69}=inp_8[17]+inp_9[16]+inp_10[15];
  assign {FA_cout_70,FA_out_70}=inp_8[20]+inp_9[19]+inp_10[18];
  assign {FA_cout_71,FA_out_71}=inp_8[23]+inp_9[22]+inp_10[21];
  assign {FA_cout_72,FA_out_72}=inp_9[2]+inp_10[1]+inp_11[0];
  assign {FA_cout_73,FA_out_73}=inp_9[3]+inp_10[2]+inp_11[1];
  assign {FA_cout_74,FA_out_74}=inp_9[4]+inp_10[3]+inp_11[2];
  assign {FA_cout_75,FA_out_75}=inp_9[5]+inp_10[4]+inp_11[3];
  assign {FA_cout_76,FA_out_76}=inp_9[6]+inp_10[5]+inp_11[4];
  assign {FA_cout_77,FA_out_77}=inp_9[7]+inp_10[6]+inp_11[5];
  assign {FA_cout_78,FA_out_78}=inp_9[8]+inp_10[7]+inp_11[6];
  assign {FA_cout_79,FA_out_79}=inp_9[9]+inp_10[8]+inp_11[7];
  assign {FA_cout_80,FA_out_80}=inp_9[10]+inp_10[9]+inp_11[8];
  assign {FA_cout_81,FA_out_81}=inp_9[11]+inp_10[10]+inp_11[9];
  assign {FA_cout_82,FA_out_82}=inp_9[12]+inp_10[11]+inp_11[10];
  assign {FA_cout_83,FA_out_83}=inp_9[13]+inp_10[12]+inp_11[11];
  assign {FA_cout_84,FA_out_84}=inp_9[14]+inp_10[13]+inp_11[12];
  assign {FA_cout_85,FA_out_85}=inp_9[17]+inp_10[16]+inp_11[15];
  assign {FA_cout_86,FA_out_86}=inp_9[20]+inp_10[19]+inp_11[18];
  assign {FA_cout_87,FA_out_87}=inp_9[23]+inp_10[22]+inp_11[21];
  assign {FA_cout_88,FA_out_88}=inp_10[14]+inp_11[13]+inp_12[12];
  assign {FA_cout_89,FA_out_89}=inp_10[17]+inp_11[16]+inp_12[15];
  assign {FA_cout_90,FA_out_90}=inp_10[20]+inp_11[19]+inp_12[18];
  assign {FA_cout_91,FA_out_91}=inp_10[23]+inp_11[22]+inp_12[21];
  assign {FA_cout_92,FA_out_92}=inp_11[14]+inp_12[13]+inp_13[12];
  assign {FA_cout_93,FA_out_93}=inp_11[17]+inp_12[16]+inp_13[15];
  assign {FA_cout_94,FA_out_94}=inp_11[20]+inp_12[19]+inp_13[18];
  assign {FA_cout_95,FA_out_95}=inp_11[23]+inp_12[22]+inp_13[21];
  assign {FA_cout_96,FA_out_96}=inp_12[2]+inp_13[1]+inp_14[0];
  assign {FA_cout_97,FA_out_97}=inp_12[3]+inp_13[2]+inp_14[1];
  assign {FA_cout_98,FA_out_98}=inp_12[4]+inp_13[3]+inp_14[2];
  assign {FA_cout_99,FA_out_99}=inp_12[5]+inp_13[4]+inp_14[3];
  assign {FA_cout_100,FA_out_100}=inp_12[6]+inp_13[5]+inp_14[4];
  assign {FA_cout_101,FA_out_101}=inp_12[7]+inp_13[6]+inp_14[5];
  assign {FA_cout_102,FA_out_102}=inp_12[8]+inp_13[7]+inp_14[6];
  assign {FA_cout_103,FA_out_103}=inp_12[9]+inp_13[8]+inp_14[7];
  assign {FA_cout_104,FA_out_104}=inp_12[10]+inp_13[9]+inp_14[8];
  assign {FA_cout_105,FA_out_105}=inp_12[11]+inp_13[10]+inp_14[9];
  assign {FA_cout_106,FA_out_106}=inp_12[14]+inp_13[13]+inp_14[12];
  assign {FA_cout_107,FA_out_107}=inp_12[17]+inp_13[16]+inp_14[15];
  assign {FA_cout_108,FA_out_108}=inp_12[20]+inp_13[19]+inp_14[18];
  assign {FA_cout_109,FA_out_109}=inp_12[23]+inp_13[22]+inp_14[21];
  assign {FA_cout_110,FA_out_110}=inp_13[11]+inp_14[10]+inp_15[9];
  assign {FA_cout_111,FA_out_111}=inp_13[14]+inp_14[13]+inp_15[12];
  assign {FA_cout_112,FA_out_112}=inp_13[17]+inp_14[16]+inp_15[15];
  assign {FA_cout_113,FA_out_113}=inp_13[20]+inp_14[19]+inp_15[18];
  assign {FA_cout_114,FA_out_114}=inp_13[23]+inp_14[22]+inp_15[21];
  assign {FA_cout_115,FA_out_115}=inp_14[11]+inp_15[10]+inp_16[9];
  assign {FA_cout_116,FA_out_116}=inp_14[14]+inp_15[13]+inp_16[12];
  assign {FA_cout_117,FA_out_117}=inp_14[17]+inp_15[16]+inp_16[15];
  assign {FA_cout_118,FA_out_118}=inp_14[20]+inp_15[19]+inp_16[18];
  assign {FA_cout_119,FA_out_119}=inp_14[23]+inp_15[22]+inp_16[21];
  assign {FA_cout_120,FA_out_120}=inp_15[2]+inp_16[1]+inp_17[0];
  assign {FA_cout_121,FA_out_121}=inp_15[3]+inp_16[2]+inp_17[1];
  assign {FA_cout_122,FA_out_122}=inp_15[4]+inp_16[3]+inp_17[2];
  assign {FA_cout_123,FA_out_123}=inp_15[5]+inp_16[4]+inp_17[3];
  assign {FA_cout_124,FA_out_124}=inp_15[6]+inp_16[5]+inp_17[4];
  assign {FA_cout_125,FA_out_125}=inp_15[7]+inp_16[6]+inp_17[5];
  assign {FA_cout_126,FA_out_126}=inp_15[8]+inp_16[7]+inp_17[6];
  assign {FA_cout_127,FA_out_127}=inp_15[11]+inp_16[10]+inp_17[9];
  assign {FA_cout_128,FA_out_128}=inp_15[14]+inp_16[13]+inp_17[12];
  assign {FA_cout_129,FA_out_129}=inp_15[17]+inp_16[16]+inp_17[15];
  assign {FA_cout_130,FA_out_130}=inp_15[20]+inp_16[19]+inp_17[18];
  assign {FA_cout_131,FA_out_131}=inp_15[23]+inp_16[22]+inp_17[21];
  assign {FA_cout_132,FA_out_132}=inp_16[8]+inp_17[7]+inp_18[6];
  assign {FA_cout_133,FA_out_133}=inp_16[11]+inp_17[10]+inp_18[9];
  assign {FA_cout_134,FA_out_134}=inp_16[14]+inp_17[13]+inp_18[12];
  assign {FA_cout_135,FA_out_135}=inp_16[17]+inp_17[16]+inp_18[15];
  assign {FA_cout_136,FA_out_136}=inp_16[20]+inp_17[19]+inp_18[18];
  assign {FA_cout_137,FA_out_137}=inp_16[23]+inp_17[22]+inp_18[21];
  assign {FA_cout_138,FA_out_138}=inp_17[8]+inp_18[7]+inp_19[6];
  assign {FA_cout_139,FA_out_139}=inp_17[11]+inp_18[10]+inp_19[9];
  assign {FA_cout_140,FA_out_140}=inp_17[14]+inp_18[13]+inp_19[12];
  assign {FA_cout_141,FA_out_141}=inp_17[17]+inp_18[16]+inp_19[15];
  assign {FA_cout_142,FA_out_142}=inp_17[20]+inp_18[19]+inp_19[18];
  assign {FA_cout_143,FA_out_143}=inp_17[23]+inp_18[22]+inp_19[21];
  assign {FA_cout_144,FA_out_144}=inp_18[2]+inp_19[1]+inp_20[0];
  assign {FA_cout_145,FA_out_145}=inp_18[3]+inp_19[2]+inp_20[1];
  assign {FA_cout_146,FA_out_146}=inp_18[4]+inp_19[3]+inp_20[2];
  assign {FA_cout_147,FA_out_147}=inp_18[5]+inp_19[4]+inp_20[3];
  assign {FA_cout_148,FA_out_148}=inp_18[8]+inp_19[7]+inp_20[6];
  assign {FA_cout_149,FA_out_149}=inp_18[11]+inp_19[10]+inp_20[9];
  assign {FA_cout_150,FA_out_150}=inp_18[14]+inp_19[13]+inp_20[12];
  assign {FA_cout_151,FA_out_151}=inp_18[17]+inp_19[16]+inp_20[15];
  assign {FA_cout_152,FA_out_152}=inp_18[20]+inp_19[19]+inp_20[18];
  assign {FA_cout_153,FA_out_153}=inp_18[23]+inp_19[22]+inp_20[21];
  assign {FA_cout_154,FA_out_154}=inp_19[5]+inp_20[4]+inp_21[3];
  assign {FA_cout_155,FA_out_155}=inp_19[8]+inp_20[7]+inp_21[6];
  assign {FA_cout_156,FA_out_156}=inp_19[11]+inp_20[10]+inp_21[9];
  assign {FA_cout_157,FA_out_157}=inp_19[14]+inp_20[13]+inp_21[12];
  assign {FA_cout_158,FA_out_158}=inp_19[17]+inp_20[16]+inp_21[15];
  assign {FA_cout_159,FA_out_159}=inp_19[20]+inp_20[19]+inp_21[18];
  assign {FA_cout_160,FA_out_160}=inp_19[23]+inp_20[22]+inp_21[21];
  assign {FA_cout_161,FA_out_161}=inp_20[5]+inp_21[4]+inp_22[3];
  assign {FA_cout_162,FA_out_162}=inp_20[8]+inp_21[7]+inp_22[6];
  assign {FA_cout_163,FA_out_163}=inp_20[11]+inp_21[10]+inp_22[9];
  assign {FA_cout_164,FA_out_164}=inp_20[14]+inp_21[13]+inp_22[12];
  assign {FA_cout_165,FA_out_165}=inp_20[17]+inp_21[16]+inp_22[15];
  assign {FA_cout_166,FA_out_166}=inp_20[20]+inp_21[19]+inp_22[18];
  assign {FA_cout_167,FA_out_167}=inp_20[23]+inp_21[22]+inp_22[21];
  assign {FA_cout_168,FA_out_168}=inp_21[2]+inp_22[1]+inp_23[0];
  assign {FA_cout_169,FA_out_169}=inp_21[5]+inp_22[4]+inp_23[3];
  assign {FA_cout_170,FA_out_170}=inp_21[8]+inp_22[7]+inp_23[6];
  assign {FA_cout_171,FA_out_171}=inp_21[11]+inp_22[10]+inp_23[9];
  assign {FA_cout_172,FA_out_172}=inp_21[14]+inp_22[13]+inp_23[12];
  assign {FA_cout_173,FA_out_173}=inp_21[17]+inp_22[16]+inp_23[15];
  assign {FA_cout_174,FA_out_174}=inp_21[20]+inp_22[19]+inp_23[18];
  assign {FA_cout_175,FA_out_175}=inp_21[23]+inp_22[22]+inp_23[21];
  assign {FA_cout_176,FA_out_176}=FA_cout_0+FA_out_1+inp_3[0];
  assign {FA_cout_177,FA_out_177}=FA_cout_1+FA_out_2+HA_out_1;
  assign {FA_cout_178,FA_out_178}=FA_cout_2+FA_out_3+HA_cout_1;
  assign {FA_cout_179,FA_out_179}=FA_cout_3+FA_out_4+FA_cout_24;
  assign {FA_cout_180,FA_out_180}=FA_cout_4+FA_out_5+FA_cout_25;
  assign {FA_cout_181,FA_out_181}=FA_cout_5+FA_out_6+FA_cout_26;
  assign {FA_cout_182,FA_out_182}=FA_cout_6+FA_out_7+FA_cout_27;
  assign {FA_cout_183,FA_out_183}=FA_cout_7+FA_out_8+FA_cout_28;
  assign {FA_cout_184,FA_out_184}=FA_cout_8+FA_out_9+FA_cout_29;
  assign {FA_cout_185,FA_out_185}=FA_cout_9+FA_out_10+FA_cout_30;
  assign {FA_cout_186,FA_out_186}=FA_cout_10+FA_out_11+FA_cout_31;
  assign {FA_cout_187,FA_out_187}=FA_cout_11+FA_out_12+FA_cout_32;
  assign {FA_cout_188,FA_out_188}=FA_cout_12+FA_out_13+FA_cout_33;
  assign {FA_cout_189,FA_out_189}=FA_cout_13+FA_out_14+FA_cout_34;
  assign {FA_cout_190,FA_out_190}=FA_cout_14+FA_out_15+FA_cout_35;
  assign {FA_cout_191,FA_out_191}=FA_cout_15+FA_out_16+FA_cout_36;
  assign {FA_cout_192,FA_out_192}=FA_cout_16+FA_out_17+FA_cout_37;
  assign {FA_cout_193,FA_out_193}=FA_cout_17+FA_out_18+FA_cout_38;
  assign {FA_cout_194,FA_out_194}=FA_cout_18+FA_out_19+FA_cout_39;
  assign {FA_cout_195,FA_out_195}=FA_cout_19+FA_out_20+FA_cout_40;
  assign {FA_cout_196,FA_out_196}=FA_cout_20+FA_out_21+FA_cout_41;
  assign {FA_cout_197,FA_out_197}=FA_cout_21+FA_out_22+FA_cout_42;
  assign {FA_cout_198,FA_out_198}=FA_cout_22+FA_out_23+FA_cout_44;
  assign {FA_cout_199,FA_out_199}=FA_cout_23+FA_out_43+FA_cout_46;
  assign {FA_cout_200,FA_out_200}=FA_cout_43+FA_out_45+FA_cout_64;
  assign {FA_cout_201,FA_out_201}=FA_out_27+HA_cout_2+FA_out_48;
  assign {FA_cout_202,FA_out_202}=FA_out_28+FA_cout_48+FA_out_49;
  assign {FA_cout_203,FA_out_203}=FA_out_29+FA_cout_49+FA_out_50;
  assign {FA_cout_204,FA_out_204}=FA_out_30+FA_cout_50+FA_out_51;
  assign {FA_cout_205,FA_out_205}=FA_out_31+FA_cout_51+FA_out_52;
  assign {FA_cout_206,FA_out_206}=FA_out_32+FA_cout_52+FA_out_53;
  assign {FA_cout_207,FA_out_207}=FA_out_33+FA_cout_53+FA_out_54;
  assign {FA_cout_208,FA_out_208}=FA_out_34+FA_cout_54+FA_out_55;
  assign {FA_cout_209,FA_out_209}=FA_out_35+FA_cout_55+FA_out_56;
  assign {FA_cout_210,FA_out_210}=FA_out_36+FA_cout_56+FA_out_57;
  assign {FA_cout_211,FA_out_211}=FA_out_37+FA_cout_57+FA_out_58;
  assign {FA_cout_212,FA_out_212}=FA_out_38+FA_cout_58+FA_out_59;
  assign {FA_cout_213,FA_out_213}=FA_out_39+FA_cout_59+FA_out_60;
  assign {FA_cout_214,FA_out_214}=FA_out_40+FA_cout_60+FA_out_61;
  assign {FA_cout_215,FA_out_215}=FA_out_41+FA_cout_61+FA_out_62;
  assign {FA_cout_216,FA_out_216}=FA_out_42+FA_cout_62+FA_out_63;
  assign {FA_cout_217,FA_out_217}=FA_out_44+FA_cout_63+FA_out_66;
  assign {FA_cout_218,FA_out_218}=FA_cout_45+FA_out_47+FA_cout_67;
  assign {FA_cout_219,FA_out_219}=FA_out_46+FA_cout_66+FA_out_69;
  assign {FA_cout_220,FA_out_220}=FA_cout_47+FA_out_65+FA_cout_70;
  assign {FA_cout_221,FA_out_221}=FA_out_64+FA_cout_69+FA_out_85;
  assign {FA_cout_222,FA_out_222}=FA_cout_65+FA_out_68+FA_cout_86;
  assign {FA_cout_223,FA_out_223}=FA_out_67+FA_cout_85+FA_out_89;
  assign {FA_cout_224,FA_out_224}=FA_cout_68+FA_out_71+FA_cout_90;
  assign {FA_cout_225,FA_out_225}=FA_out_70+FA_cout_89+FA_out_93;
  assign {FA_cout_226,FA_out_226}=FA_cout_71+FA_out_87+FA_cout_94;
  assign {FA_cout_227,FA_out_227}=FA_cout_72+FA_out_73+inp_12[0];
  assign {FA_cout_228,FA_out_228}=FA_cout_73+FA_out_74+HA_out_4;
  assign {FA_cout_229,FA_out_229}=FA_cout_74+FA_out_75+HA_cout_4;
  assign {FA_cout_230,FA_out_230}=FA_cout_75+FA_out_76+FA_cout_96;
  assign {FA_cout_231,FA_out_231}=FA_cout_76+FA_out_77+FA_cout_97;
  assign {FA_cout_232,FA_out_232}=FA_cout_77+FA_out_78+FA_cout_98;
  assign {FA_cout_233,FA_out_233}=FA_cout_78+FA_out_79+FA_cout_99;
  assign {FA_cout_234,FA_out_234}=FA_cout_79+FA_out_80+FA_cout_100;
  assign {FA_cout_235,FA_out_235}=FA_cout_80+FA_out_81+FA_cout_101;
  assign {FA_cout_236,FA_out_236}=FA_cout_81+FA_out_82+FA_cout_102;
  assign {FA_cout_237,FA_out_237}=FA_cout_82+FA_out_83+FA_cout_103;
  assign {FA_cout_238,FA_out_238}=FA_cout_83+FA_out_84+FA_cout_104;
  assign {FA_cout_239,FA_out_239}=FA_cout_84+FA_out_88+FA_cout_105;
  assign {FA_cout_240,FA_out_240}=FA_out_86+FA_cout_93+FA_out_107;
  assign {FA_cout_241,FA_out_241}=FA_cout_87+FA_out_91+FA_cout_108;
  assign {FA_cout_242,FA_out_242}=FA_cout_88+FA_out_92+FA_cout_110;
  assign {FA_cout_243,FA_out_243}=FA_out_90+FA_cout_107+FA_out_112;
  assign {FA_cout_244,FA_out_244}=FA_cout_91+FA_out_95+FA_cout_113;
  assign {FA_cout_245,FA_out_245}=FA_cout_92+FA_out_106+FA_cout_115;
  assign {FA_cout_246,FA_out_246}=FA_out_94+FA_cout_112+FA_out_117;
  assign {FA_cout_247,FA_out_247}=FA_cout_95+FA_out_109+FA_cout_118;
  assign {FA_cout_248,FA_out_248}=FA_cout_106+FA_out_111+FA_cout_127;
  assign {FA_cout_249,FA_out_249}=FA_out_108+FA_cout_117+FA_out_129;
  assign {FA_cout_250,FA_out_250}=FA_cout_109+FA_out_114+FA_cout_130;
  assign {FA_cout_251,FA_out_251}=FA_out_99+HA_cout_5+FA_out_120;
  assign {FA_cout_252,FA_out_252}=FA_out_100+FA_cout_120+FA_out_121;
  assign {FA_cout_253,FA_out_253}=FA_out_101+FA_cout_121+FA_out_122;
  assign {FA_cout_254,FA_out_254}=FA_out_102+FA_cout_122+FA_out_123;
  assign {FA_cout_255,FA_out_255}=FA_out_103+FA_cout_123+FA_out_124;
  assign {FA_cout_256,FA_out_256}=FA_out_104+FA_cout_124+FA_out_125;
  assign {FA_cout_257,FA_out_257}=FA_out_105+FA_cout_125+FA_out_126;
  assign {FA_cout_258,FA_out_258}=FA_out_110+FA_cout_126+FA_out_132;
  assign {FA_cout_259,FA_out_259}=FA_cout_111+FA_out_116+FA_cout_133;
  assign {FA_cout_260,FA_out_260}=FA_out_113+FA_cout_129+FA_out_135;
  assign {FA_cout_261,FA_out_261}=FA_cout_114+FA_out_119+FA_cout_136;
  assign {FA_cout_262,FA_out_262}=FA_out_115+FA_cout_132+FA_out_138;
  assign {FA_cout_263,FA_out_263}=FA_cout_116+FA_out_128+FA_cout_139;
  assign {FA_cout_264,FA_out_264}=FA_out_118+FA_cout_135+FA_out_141;
  assign {FA_cout_265,FA_out_265}=FA_cout_119+FA_out_131+FA_cout_142;
  assign {FA_cout_266,FA_out_266}=FA_out_127+FA_cout_138+FA_out_148;
  assign {FA_cout_267,FA_out_267}=FA_cout_128+FA_out_134+FA_cout_149;
  assign {FA_cout_268,FA_out_268}=FA_out_130+FA_cout_141+FA_out_151;
  assign {FA_cout_269,FA_out_269}=FA_cout_131+FA_out_137+FA_cout_152;
  assign {FA_cout_270,FA_out_270}=FA_out_133+FA_cout_148+FA_out_155;
  assign {FA_cout_271,FA_out_271}=FA_cout_134+FA_out_140+FA_cout_156;
  assign {FA_cout_272,FA_out_272}=FA_out_136+FA_cout_151+FA_out_158;
  assign {FA_cout_273,FA_out_273}=FA_cout_137+FA_out_143+FA_cout_159;
  assign {FA_cout_274,FA_out_274}=FA_out_139+FA_cout_155+FA_out_162;
  assign {FA_cout_275,FA_out_275}=FA_cout_140+FA_out_150+FA_cout_163;
  assign {FA_cout_276,FA_out_276}=FA_out_142+FA_cout_158+FA_out_165;
  assign {FA_cout_277,FA_out_277}=FA_cout_143+FA_out_153+FA_cout_166;
  assign {FA_cout_278,FA_out_278}=FA_cout_144+FA_out_145+inp_21[0];
  assign {FA_cout_279,FA_out_279}=FA_cout_145+FA_out_146+HA_out_7;
  assign {FA_cout_280,FA_out_280}=FA_cout_146+FA_out_147+HA_cout_7;
  assign {FA_cout_281,FA_out_281}=FA_cout_147+FA_out_154+FA_cout_168;
  assign {FA_cout_282,FA_out_282}=FA_out_149+FA_cout_162+FA_out_170;
  assign {FA_cout_283,FA_out_283}=FA_cout_150+FA_out_157+FA_cout_171;
  assign {FA_cout_284,FA_out_284}=FA_out_152+FA_cout_165+FA_out_173;
  assign {FA_cout_285,FA_out_285}=FA_cout_153+FA_out_160+FA_cout_174;
  assign {FA_cout_286,FA_out_286}=FA_cout_154+FA_out_161+HA_cout_8;
  assign {FA_cout_287,FA_out_287}=FA_out_156+FA_cout_170+HA_out_10;
  assign {FA_cout_288,FA_out_288}=FA_cout_157+FA_out_164+HA_cout_11;
  assign {FA_cout_289,FA_out_289}=FA_out_159+FA_cout_173+HA_out_13;
  assign {FA_cout_290,FA_out_290}=FA_cout_160+FA_out_167+HA_cout_14;
  assign {FA_cout_291,FA_out_291}=FA_out_163+HA_cout_10+inp_23[8];
  assign {FA_cout_292,FA_out_292}=FA_out_166+HA_cout_13+inp_23[17];
  assign {FA_cout_293,FA_out_293}=REGS_5+REGS_28+REGS_54;
  assign {FA_cout_294,FA_out_294}=REGS_6+REGS_29+REGS_55;
  assign {FA_cout_295,FA_out_295}=REGS_7+REGS_30+REGS_56;
  assign {FA_cout_296,FA_out_296}=REGS_8+REGS_31+REGS_57;
  assign {FA_cout_297,FA_out_297}=REGS_9+REGS_32+REGS_58;
  assign {FA_cout_298,FA_out_298}=REGS_10+REGS_33+REGS_59;
  assign {FA_cout_299,FA_out_299}=REGS_11+REGS_34+REGS_60;
  assign {FA_cout_300,FA_out_300}=REGS_12+REGS_35+REGS_61;
  assign {FA_cout_301,FA_out_301}=REGS_13+REGS_36+REGS_62;
  assign {FA_cout_302,FA_out_302}=REGS_14+REGS_37+REGS_63;
  assign {FA_cout_303,FA_out_303}=REGS_15+REGS_38+REGS_64;
  assign {FA_cout_304,FA_out_304}=REGS_16+REGS_39+REGS_65;
  assign {FA_cout_305,FA_out_305}=REGS_17+REGS_40+REGS_66;
  assign {FA_cout_306,FA_out_306}=REGS_18+REGS_41+REGS_67;
  assign {FA_cout_307,FA_out_307}=REGS_19+REGS_42+REGS_68;
  assign {FA_cout_308,FA_out_308}=REGS_20+REGS_43+REGS_69;
  assign {FA_cout_309,FA_out_309}=REGS_21+REGS_44+REGS_70;
  assign {FA_cout_310,FA_out_310}=REGS_22+REGS_45+REGS_71;
  assign {FA_cout_311,FA_out_311}=REGS_23+REGS_46+REGS_72;
  assign {FA_cout_312,FA_out_312}=REGS_24+REGS_47+REGS_73;
  assign {FA_cout_313,FA_out_313}=REGS_25+REGS_48+REGS_74;
  assign {FA_cout_314,FA_out_314}=REGS_49+REGS_50+REGS_96;
  assign {FA_cout_315,FA_out_315}=REGS_51+REGS_52+REGS_100;
  assign {FA_cout_316,FA_out_316}=REGS_53+REGS_75+REGS_104;
  assign {FA_cout_317,FA_out_317}=REGS_76+REGS_97+REGS_108;
  assign {FA_cout_318,FA_out_318}=REGS_82+REGS_114+REGS_132;
  assign {FA_cout_319,FA_out_319}=REGS_83+REGS_115+REGS_133;
  assign {FA_cout_320,FA_out_320}=REGS_84+REGS_116+REGS_134;
  assign {FA_cout_321,FA_out_321}=REGS_85+REGS_117+REGS_135;
  assign {FA_cout_322,FA_out_322}=REGS_86+REGS_118+REGS_136;
  assign {FA_cout_323,FA_out_323}=REGS_87+REGS_119+REGS_137;
  assign {FA_cout_324,FA_out_324}=REGS_88+REGS_120+REGS_138;
  assign {FA_cout_325,FA_out_325}=REGS_89+REGS_121+REGS_139;
  assign {FA_cout_326,FA_out_326}=REGS_90+REGS_122+REGS_140;
  assign {FA_cout_327,FA_out_327}=REGS_91+REGS_123+REGS_141;
  assign {FA_cout_328,FA_out_328}=REGS_92+REGS_124+REGS_142;
  assign {FA_cout_329,FA_out_329}=REGS_93+REGS_125+REGS_143;
  assign {FA_cout_330,FA_out_330}=REGS_94+REGS_126+REGS_144;
  assign {FA_cout_331,FA_out_331}=REGS_95+REGS_127+REGS_145;
  assign {FA_cout_332,FA_out_332}=REGS_98+REGS_101+REGS_129;
  assign {FA_cout_333,FA_out_333}=REGS_99+REGS_146+REGS_151;
  assign {FA_cout_334,FA_out_334}=REGS_102+REGS_105+REGS_148;
  assign {FA_cout_335,FA_out_335}=REGS_103+REGS_152+REGS_157;
  assign {FA_cout_336,FA_out_336}=REGS_106+REGS_109+REGS_154;
  assign {FA_cout_337,FA_out_337}=REGS_107+REGS_158+REGS_175;
  assign {FA_cout_338,FA_out_338}=REGS_110+REGS_130+REGS_160;
  assign {FA_cout_339,FA_out_339}=REGS_128+REGS_176+REGS_192;
  assign {FA_cout_340,FA_out_340}=REGS_131+REGS_149+REGS_178;
  assign {FA_cout_341,FA_out_341}=REGS_147+REGS_193+REGS_200;
  assign {FA_cout_342,FA_out_342}=REGS_150+REGS_155+REGS_195;
  assign {FA_cout_343,FA_out_343}=REGS_153+REGS_201+REGS_208;
  assign {FA_cout_344,FA_out_344}=REGS_156+REGS_161+REGS_203;
  assign {FA_cout_345,FA_out_345}=REGS_159+REGS_209+REGS_216;
  assign {FA_cout_346,FA_out_346}=REGS_162+REGS_179+REGS_211;
  assign {FA_cout_347,FA_out_347}=REGS_167+REGS_183+REGS_222;
  assign {FA_cout_348,FA_out_348}=REGS_168+REGS_184+REGS_223;
  assign {FA_cout_349,FA_out_349}=REGS_169+REGS_185+REGS_224;
  assign {FA_cout_350,FA_out_350}=REGS_170+REGS_186+REGS_225;
  assign {FA_cout_351,FA_out_351}=REGS_171+REGS_187+REGS_226;
  assign {FA_cout_352,FA_out_352}=REGS_172+REGS_188+REGS_227;
  assign {FA_cout_353,FA_out_353}=REGS_173+REGS_189+REGS_228;
  assign {FA_cout_354,FA_out_354}=REGS_174+REGS_190+REGS_229;
  assign {FA_cout_355,FA_out_355}=REGS_177+REGS_217+REGS_232;
  assign {FA_cout_356,FA_out_356}=REGS_180+REGS_196+REGS_219;
  assign {FA_cout_357,FA_out_357}=REGS_191+REGS_198+REGS_243;
  assign {FA_cout_358,FA_out_358}=REGS_194+REGS_233+REGS_246;
  assign {FA_cout_359,FA_out_359}=REGS_197+REGS_204+REGS_235;
  assign {FA_cout_360,FA_out_360}=REGS_199+REGS_206+REGS_253;
  assign {FA_cout_361,FA_out_361}=REGS_202+REGS_247+REGS_256;
  assign {FA_cout_362,FA_out_362}=REGS_205+REGS_212+REGS_249;
  assign {FA_cout_363,FA_out_363}=REGS_207+REGS_214+REGS_263;
  assign {FA_cout_364,FA_out_364}=REGS_210+REGS_257+REGS_265;
  assign {FA_cout_365,FA_out_365}=REGS_213+REGS_220+REGS_259;
  assign {FA_cout_366,FA_out_366}=REGS_215+REGS_230+REGS_273;
  assign {FA_cout_367,FA_out_367}=REGS_218+REGS_266+REGS_275;
  assign {FA_cout_368,FA_out_368}=REGS_221+REGS_236+REGS_277;
  assign {FA_cout_369,FA_out_369}=REGS_237+REGS_250+REGS_282;
  assign {FA_cout_370,FA_out_370}=FA_cout_294+FA_out_295+REGS_77;
  assign {FA_cout_371,FA_out_371}=FA_cout_295+FA_out_296+REGS_78;
  assign {FA_cout_372,FA_out_372}=FA_cout_296+FA_out_297+HA_out_34;
  assign {FA_cout_373,FA_out_373}=FA_cout_297+FA_out_298+HA_cout_34;
  assign {FA_cout_374,FA_out_374}=FA_cout_298+FA_out_299+HA_cout_35;
  assign {FA_cout_375,FA_out_375}=FA_cout_299+FA_out_300+HA_cout_36;
  assign {FA_cout_376,FA_out_376}=FA_cout_300+FA_out_301+FA_cout_318;
  assign {FA_cout_377,FA_out_377}=FA_cout_301+FA_out_302+FA_cout_319;
  assign {FA_cout_378,FA_out_378}=FA_cout_302+FA_out_303+FA_cout_320;
  assign {FA_cout_379,FA_out_379}=FA_cout_303+FA_out_304+FA_cout_321;
  assign {FA_cout_380,FA_out_380}=FA_cout_304+FA_out_305+FA_cout_322;
  assign {FA_cout_381,FA_out_381}=FA_cout_305+FA_out_306+FA_cout_323;
  assign {FA_cout_382,FA_out_382}=FA_cout_306+FA_out_307+FA_cout_324;
  assign {FA_cout_383,FA_out_383}=FA_cout_307+FA_out_308+FA_cout_325;
  assign {FA_cout_384,FA_out_384}=FA_cout_308+FA_out_309+FA_cout_326;
  assign {FA_cout_385,FA_out_385}=FA_cout_309+FA_out_310+FA_cout_327;
  assign {FA_cout_386,FA_out_386}=FA_cout_310+FA_out_311+FA_cout_328;
  assign {FA_cout_387,FA_out_387}=FA_cout_311+FA_out_312+FA_cout_329;
  assign {FA_cout_388,FA_out_388}=FA_cout_312+FA_out_313+FA_cout_330;
  assign {FA_cout_389,FA_out_389}=FA_cout_313+FA_out_314+FA_cout_331;
  assign {FA_cout_390,FA_out_390}=FA_cout_314+FA_out_315+FA_cout_333;
  assign {FA_cout_391,FA_out_391}=FA_cout_315+FA_out_316+FA_cout_335;
  assign {FA_cout_392,FA_out_392}=FA_cout_316+FA_out_317+FA_cout_337;
  assign {FA_cout_393,FA_out_393}=FA_cout_317+FA_out_332+FA_cout_339;
  assign {FA_cout_394,FA_out_394}=FA_cout_332+FA_out_334+FA_cout_341;
  assign {FA_cout_395,FA_out_395}=FA_out_323+HA_cout_37+HA_out_38;
  assign {FA_cout_396,FA_out_396}=FA_out_324+HA_cout_38+FA_out_347;
  assign {FA_cout_397,FA_out_397}=FA_out_325+FA_cout_347+FA_out_348;
  assign {FA_cout_398,FA_out_398}=FA_out_326+FA_cout_348+FA_out_349;
  assign {FA_cout_399,FA_out_399}=FA_out_327+FA_cout_349+FA_out_350;
  assign {FA_cout_400,FA_out_400}=FA_out_328+FA_cout_350+FA_out_351;
  assign {FA_cout_401,FA_out_401}=FA_out_329+FA_cout_351+FA_out_352;
  assign {FA_cout_402,FA_out_402}=FA_out_330+FA_cout_352+FA_out_353;
  assign {FA_cout_403,FA_out_403}=FA_out_331+FA_cout_353+FA_out_354;
  assign {FA_cout_404,FA_out_404}=FA_out_333+FA_cout_354+FA_out_357;
  assign {FA_cout_405,FA_out_405}=FA_cout_334+FA_out_336+FA_cout_343;
  assign {FA_cout_406,FA_out_406}=FA_out_335+FA_cout_357+FA_out_360;
  assign {FA_cout_407,FA_out_407}=FA_cout_336+FA_out_338+FA_cout_345;
  assign {FA_cout_408,FA_out_408}=FA_out_337+FA_cout_360+FA_out_363;
  assign {FA_cout_409,FA_out_409}=FA_cout_338+FA_out_340+FA_cout_355;
  assign {FA_cout_410,FA_out_410}=FA_out_339+FA_cout_363+FA_out_366;
  assign {FA_cout_411,FA_out_411}=FA_cout_340+FA_out_342+FA_cout_358;
  assign {FA_cout_412,FA_out_412}=FA_out_341+FA_cout_366+HA_out_39;
  assign {FA_cout_413,FA_out_413}=FA_cout_342+FA_out_344+FA_cout_361;
  assign {FA_cout_414,FA_out_414}=FA_out_343+HA_cout_39+HA_out_44;
  assign {FA_cout_415,FA_out_415}=FA_cout_344+FA_out_346+FA_cout_364;
  assign {FA_cout_416,FA_out_416}=FA_out_345+HA_cout_44+HA_out_46;
  assign {FA_cout_417,FA_out_417}=FA_cout_346+FA_out_356+FA_cout_367;
  assign {FA_cout_418,FA_out_418}=FA_out_355+HA_cout_46+REGS_274;
  assign {FA_cout_419,FA_out_419}=FA_cout_356+FA_out_359+HA_cout_40;
  assign {FA_cout_420,FA_out_420}=FA_cout_359+FA_out_362+REGS_258;
  assign {FA_cout_421,FA_out_421}=FA_cout_362+FA_out_365+REGS_267;
  assign {FA_cout_422,FA_out_422}=FA_cout_372+FA_out_373+HA_out_35;
  assign {FA_cout_423,FA_out_423}=FA_cout_373+FA_out_374+HA_out_36;
  assign {FA_cout_424,FA_out_424}=FA_cout_374+FA_out_375+FA_out_318;
  assign {FA_cout_425,FA_out_425}=FA_cout_375+FA_out_376+FA_out_319;
  assign {FA_cout_426,FA_out_426}=FA_cout_376+FA_out_377+HA_out_52;
  assign {FA_cout_427,FA_out_427}=FA_cout_377+FA_out_378+HA_cout_52;
  assign {FA_cout_428,FA_out_428}=FA_cout_378+FA_out_379+HA_cout_53;
  assign {FA_cout_429,FA_out_429}=FA_cout_379+FA_out_380+HA_cout_54;
  assign {FA_cout_430,FA_out_430}=FA_cout_380+FA_out_381+FA_cout_395;
  assign {FA_cout_431,FA_out_431}=FA_cout_381+FA_out_382+FA_cout_396;
  assign {FA_cout_432,FA_out_432}=FA_cout_382+FA_out_383+FA_cout_397;
  assign {FA_cout_433,FA_out_433}=FA_cout_383+FA_out_384+FA_cout_398;
  assign {FA_cout_434,FA_out_434}=FA_cout_384+FA_out_385+FA_cout_399;
  assign {FA_cout_435,FA_out_435}=FA_cout_385+FA_out_386+FA_cout_400;
  assign {FA_cout_436,FA_out_436}=FA_cout_386+FA_out_387+FA_cout_401;
  assign {FA_cout_437,FA_out_437}=FA_cout_387+FA_out_388+FA_cout_402;
  assign {FA_cout_438,FA_out_438}=FA_cout_388+FA_out_389+FA_cout_403;
  assign {FA_cout_439,FA_out_439}=FA_cout_389+FA_out_390+FA_cout_404;
  assign {FA_cout_440,FA_out_440}=FA_cout_390+FA_out_391+FA_cout_406;
  assign {FA_cout_441,FA_out_441}=FA_cout_391+FA_out_392+FA_cout_408;
  assign {FA_cout_442,FA_out_442}=FA_cout_392+FA_out_393+FA_cout_410;
  assign {FA_cout_443,FA_out_443}=FA_cout_393+FA_out_394+FA_cout_412;
  assign {FA_cout_444,FA_out_444}=FA_cout_394+FA_out_405+FA_cout_414;
  assign {FA_cout_445,FA_out_445}=FA_cout_405+FA_out_407+FA_cout_416;
  assign {FA_cout_446,FA_out_446}=FA_out_403+HA_cout_59+HA_out_60;
  assign {FA_cout_447,FA_out_447}=FA_out_404+HA_cout_60+HA_out_61;
  assign {FA_cout_448,FA_out_448}=FA_out_406+HA_cout_61+REGS_262;
  assign {FA_cout_449,FA_out_449}=FA_cout_407+FA_out_409+FA_cout_418;
  assign {FA_cout_450,FA_out_450}=FA_cout_409+FA_out_411+HA_cout_55;
  assign {FA_cout_451,FA_out_451}=FA_cout_411+FA_out_413+FA_out_364;
  assign {FA_cout_452,FA_out_452}=FA_cout_413+FA_out_415+FA_out_367;
  assign {FA_cout_453,FA_out_453}=FA_cout_415+FA_out_417+HA_out_40;
  assign {FA_cout_454,FA_out_454}=FA_cout_417+FA_out_419+REGS_248;
  assign {FA_cout_455,FA_out_455}=FA_cout_426+FA_out_427+HA_out_53;
  assign {FA_cout_456,FA_out_456}=FA_cout_427+FA_out_428+HA_out_54;
  assign {FA_cout_457,FA_out_457}=FA_cout_428+FA_out_429+FA_out_395;
  assign {FA_cout_458,FA_out_458}=FA_cout_429+FA_out_430+FA_out_396;
  assign {FA_cout_459,FA_out_459}=FA_cout_430+FA_out_431+FA_out_397;
  assign {FA_cout_460,FA_out_460}=FA_cout_431+FA_out_432+FA_out_398;
  assign {FA_cout_461,FA_out_461}=FA_cout_432+FA_out_433+HA_out_70;
  assign {FA_cout_462,FA_out_462}=FA_cout_433+FA_out_434+HA_cout_70;
  assign {FA_cout_463,FA_out_463}=FA_cout_434+FA_out_435+HA_cout_71;
  assign {FA_cout_464,FA_out_464}=FA_cout_435+FA_out_436+HA_cout_72;
  assign {FA_cout_465,FA_out_465}=FA_cout_436+FA_out_437+HA_cout_73;
  assign {FA_cout_466,FA_out_466}=FA_cout_437+FA_out_438+FA_cout_446;
  assign {FA_cout_467,FA_out_467}=FA_cout_438+FA_out_439+FA_cout_447;
  assign {FA_cout_468,FA_out_468}=FA_cout_439+FA_out_440+FA_cout_448;
  assign {FA_cout_469,FA_out_469}=FA_cout_440+FA_out_441+HA_cout_74;
  assign {FA_cout_470,FA_out_470}=FA_cout_441+FA_out_442+FA_out_412;
  assign {FA_cout_471,FA_out_471}=FA_cout_442+FA_out_443+FA_out_414;
  assign {FA_cout_472,FA_out_472}=FA_cout_443+FA_out_444+FA_out_416;
  assign {FA_cout_473,FA_out_473}=FA_cout_444+FA_out_445+FA_out_418;
  assign {FA_cout_474,FA_out_474}=FA_cout_445+FA_out_449+HA_out_55;
  assign {FA_cout_475,FA_out_475}=FA_cout_449+FA_out_450+FA_out_361;
  assign {FA_cout_476,FA_out_476}=REGS_305+REGS_328+REGS_349;
  assign {FA_cout_477,FA_out_477}=REGS_306+REGS_329+REGS_350;
  assign {FA_cout_478,FA_out_478}=REGS_307+REGS_330+REGS_351;
  assign {FA_cout_479,FA_out_479}=REGS_308+REGS_331+REGS_352;
  assign {FA_cout_480,FA_out_480}=REGS_309+REGS_332+REGS_353;
  assign {FA_cout_481,FA_out_481}=REGS_310+REGS_333+REGS_354;
  assign {FA_cout_482,FA_out_482}=REGS_311+REGS_334+REGS_355;
  assign {FA_cout_483,FA_out_483}=REGS_312+REGS_335+REGS_358;
  assign {HA_cout_0,HA_out_0}=inp_0[1]+inp_1[0];
  assign {HA_cout_1,HA_out_1}=inp_3[1]+inp_4[0];
  assign {HA_cout_2,HA_out_2}=inp_6[1]+inp_7[0];
  assign {HA_cout_3,HA_out_3}=inp_9[1]+inp_10[0];
  assign {HA_cout_4,HA_out_4}=inp_12[1]+inp_13[0];
  assign {HA_cout_5,HA_out_5}=inp_15[1]+inp_16[0];
  assign {HA_cout_6,HA_out_6}=inp_18[1]+inp_19[0];
  assign {HA_cout_7,HA_out_7}=inp_21[1]+inp_22[0];
  assign {HA_cout_8,HA_out_8}=inp_22[2]+inp_23[1];
  assign {HA_cout_9,HA_out_9}=inp_22[5]+inp_23[4];
  assign {HA_cout_10,HA_out_10}=inp_22[8]+inp_23[7];
  assign {HA_cout_11,HA_out_11}=inp_22[11]+inp_23[10];
  assign {HA_cout_12,HA_out_12}=inp_22[14]+inp_23[13];
  assign {HA_cout_13,HA_out_13}=inp_22[17]+inp_23[16];
  assign {HA_cout_14,HA_out_14}=inp_22[20]+inp_23[19];
  assign {HA_cout_15,HA_out_15}=inp_22[23]+inp_23[22];
  assign {HA_cout_16,HA_out_16}=HA_cout_0+FA_out_0;
  assign {HA_cout_17,HA_out_17}=FA_out_25+inp_6[0];
  assign {HA_cout_18,HA_out_18}=FA_out_26+HA_out_2;
  assign {HA_cout_19,HA_out_19}=HA_cout_3+FA_out_72;
  assign {HA_cout_20,HA_out_20}=FA_out_97+inp_15[0];
  assign {HA_cout_21,HA_out_21}=FA_out_98+HA_out_5;
  assign {HA_cout_22,HA_out_22}=HA_cout_6+FA_out_144;
  assign {HA_cout_23,HA_out_23}=FA_cout_161+FA_out_169;
  assign {HA_cout_24,HA_out_24}=FA_cout_164+FA_out_172;
  assign {HA_cout_25,HA_out_25}=FA_cout_167+FA_out_175;
  assign {HA_cout_26,HA_out_26}=FA_cout_169+HA_out_9;
  assign {HA_cout_27,HA_out_27}=FA_cout_172+HA_out_12;
  assign {HA_cout_28,HA_out_28}=FA_cout_175+HA_out_15;
  assign {HA_cout_29,HA_out_29}=HA_cout_9+inp_23[5];
  assign {HA_cout_30,HA_out_30}=HA_cout_12+inp_23[14];
  assign {HA_cout_31,HA_out_31}=HA_cout_15+inp_23[23];
  assign {HA_cout_32,HA_out_32}=REGS_3+REGS_26;
  assign {HA_cout_33,HA_out_33}=REGS_4+REGS_27;
  assign {HA_cout_34,HA_out_34}=REGS_79+REGS_111;
  assign {HA_cout_35,HA_out_35}=REGS_80+REGS_112;
  assign {HA_cout_36,HA_out_36}=REGS_81+REGS_113;
  assign {HA_cout_37,HA_out_37}=REGS_165+REGS_181;
  assign {HA_cout_38,HA_out_38}=REGS_166+REGS_182;
  assign {HA_cout_39,HA_out_39}=REGS_231+REGS_244;
  assign {HA_cout_40,HA_out_40}=REGS_234+REGS_276;
  assign {HA_cout_41,HA_out_41}=REGS_240+REGS_270;
  assign {HA_cout_42,HA_out_42}=REGS_241+REGS_271;
  assign {HA_cout_43,HA_out_43}=REGS_242+REGS_280;
  assign {HA_cout_44,HA_out_44}=REGS_245+REGS_254;
  assign {HA_cout_45,HA_out_45}=REGS_251+REGS_260;
  assign {HA_cout_46,HA_out_46}=REGS_255+REGS_264;
  assign {HA_cout_47,HA_out_47}=REGS_261+REGS_268;
  assign {HA_cout_48,HA_out_48}=REGS_269+REGS_278;
  assign {HA_cout_49,HA_out_49}=HA_cout_32+HA_out_33;
  assign {HA_cout_50,HA_out_50}=HA_cout_33+FA_out_293;
  assign {HA_cout_51,HA_out_51}=FA_cout_293+FA_out_294;
  assign {HA_cout_52,HA_out_52}=FA_out_320+REGS_163;
  assign {HA_cout_53,HA_out_53}=FA_out_321+REGS_164;
  assign {HA_cout_54,HA_out_54}=FA_out_322+HA_out_37;
  assign {HA_cout_55,HA_out_55}=FA_out_358+REGS_281;
  assign {HA_cout_56,HA_out_56}=FA_cout_365+FA_out_368;
  assign {HA_cout_57,HA_out_57}=FA_cout_368+FA_out_369;
  assign {HA_cout_58,HA_out_58}=FA_cout_369+HA_out_45;
  assign {HA_cout_59,HA_out_59}=HA_cout_41+HA_out_42;
  assign {HA_cout_60,HA_out_60}=HA_cout_42+HA_out_43;
  assign {HA_cout_61,HA_out_61}=HA_cout_43+REGS_252;
  assign {HA_cout_62,HA_out_62}=HA_cout_45+HA_out_47;
  assign {HA_cout_63,HA_out_63}=HA_cout_47+HA_out_48;
  assign {HA_cout_64,HA_out_64}=HA_cout_48+REGS_279;
  assign {HA_cout_65,HA_out_65}=HA_cout_49+HA_out_50;
  assign {HA_cout_66,HA_out_66}=HA_cout_50+HA_out_51;
  assign {HA_cout_67,HA_out_67}=HA_cout_51+FA_out_370;
  assign {HA_cout_68,HA_out_68}=FA_cout_370+FA_out_371;
  assign {HA_cout_69,HA_out_69}=FA_cout_371+FA_out_372;
  assign {HA_cout_70,HA_out_70}=FA_out_399+REGS_238;
  assign {HA_cout_71,HA_out_71}=FA_out_400+REGS_239;
  assign {HA_cout_72,HA_out_72}=FA_out_401+HA_out_41;
  assign {HA_cout_73,HA_out_73}=FA_out_402+HA_out_59;
  assign {HA_cout_74,HA_out_74}=FA_out_408+REGS_272;
  assign {HA_cout_75,HA_out_75}=FA_cout_419+FA_out_420;
  assign {HA_cout_76,HA_out_76}=FA_cout_420+FA_out_421;
  assign {HA_cout_77,HA_out_77}=FA_cout_421+HA_out_56;
  assign {HA_cout_78,HA_out_78}=HA_cout_56+HA_out_57;
  assign {HA_cout_79,HA_out_79}=HA_cout_57+HA_out_58;
  assign {HA_cout_80,HA_out_80}=HA_cout_58+HA_out_62;
  assign {HA_cout_81,HA_out_81}=HA_cout_62+HA_out_63;
  assign {HA_cout_82,HA_out_82}=HA_cout_63+HA_out_64;
  assign {HA_cout_83,HA_out_83}=HA_cout_65+HA_out_66;
  assign {HA_cout_84,HA_out_84}=HA_cout_66+HA_out_67;
  assign {HA_cout_85,HA_out_85}=HA_cout_67+HA_out_68;
  assign {HA_cout_86,HA_out_86}=HA_cout_68+HA_out_69;
  assign {HA_cout_87,HA_out_87}=HA_cout_69+FA_out_422;
  assign {HA_cout_88,HA_out_88}=FA_cout_422+FA_out_423;
  assign {HA_cout_89,HA_out_89}=FA_cout_423+FA_out_424;
  assign {HA_cout_90,HA_out_90}=FA_cout_424+FA_out_425;
  assign {HA_cout_91,HA_out_91}=FA_cout_425+FA_out_426;
  assign {HA_cout_92,HA_out_92}=FA_cout_450+FA_out_451;
  assign {HA_cout_93,HA_out_93}=FA_cout_451+FA_out_452;
  assign {HA_cout_94,HA_out_94}=FA_cout_452+FA_out_453;
  assign {HA_cout_95,HA_out_95}=FA_cout_453+FA_out_454;
  assign {HA_cout_96,HA_out_96}=FA_cout_454+HA_out_75;
  assign {HA_cout_97,HA_out_97}=HA_cout_75+HA_out_76;
  assign {HA_cout_98,HA_out_98}=HA_cout_76+HA_out_77;
  assign {HA_cout_99,HA_out_99}=HA_cout_77+HA_out_78;
  assign {HA_cout_100,HA_out_100}=HA_cout_78+HA_out_79;
  assign {HA_cout_101,HA_out_101}=HA_cout_79+HA_out_80;
  assign {HA_cout_102,HA_out_102}=HA_cout_80+HA_out_81;
  assign {HA_cout_103,HA_out_103}=HA_cout_81+HA_out_82;
  assign {HA_cout_104,HA_out_104}=HA_cout_82+HA_cout_64;
  assign {HA_cout_105,HA_out_105}=REGS_290+REGS_313;
  assign {HA_cout_106,HA_out_106}=REGS_291+REGS_314;
  assign {HA_cout_107,HA_out_107}=REGS_292+REGS_315;
  assign {HA_cout_108,HA_out_108}=REGS_293+REGS_316;
  assign {HA_cout_109,HA_out_109}=REGS_294+REGS_317;
  assign {HA_cout_110,HA_out_110}=REGS_295+REGS_318;
  assign {HA_cout_111,HA_out_111}=REGS_296+REGS_319;
  assign {HA_cout_112,HA_out_112}=REGS_297+REGS_320;
  assign {HA_cout_113,HA_out_113}=REGS_298+REGS_321;
  assign {HA_cout_114,HA_out_114}=REGS_299+REGS_322;
  assign {HA_cout_115,HA_out_115}=REGS_300+REGS_323;
  assign {HA_cout_116,HA_out_116}=REGS_301+REGS_324;
  assign {HA_cout_117,HA_out_117}=REGS_302+REGS_325;
  assign {HA_cout_118,HA_out_118}=REGS_303+REGS_326;
  assign {HA_cout_119,HA_out_119}=REGS_304+REGS_327;
  assign {HA_cout_120,HA_out_120}=REGS_336+REGS_337;
  assign {HA_cout_121,HA_out_121}=REGS_338+REGS_339;
  assign {HA_cout_122,HA_out_122}=REGS_340+REGS_341;
  assign {HA_cout_123,HA_out_123}=REGS_342+REGS_343;
  assign {HA_cout_124,HA_out_124}=REGS_344+REGS_345;
  assign {HA_cout_125,HA_out_125}=REGS_346+REGS_347;
  assign {HA_cout_126,HA_out_126}=REGS_348+REGS_356;
  assign {HA_cout_127,HA_out_127}=REGS_357+REGS_359;
  assign {HA_cout_128,HA_out_128}=REGS_360+REGS_361;
  assign {HA_cout_129,HA_out_129}=REGS_362+REGS_363;
  assign {HA_cout_130,HA_out_130}=REGS_364+REGS_365;
  assign {HA_cout_131,HA_out_131}=REGS_366+REGS_367;
  assign {HA_cout_132,HA_out_132}=REGS_368+REGS_369;
  assign {HA_cout_133,HA_out_133}=REGS_370+REGS_371;
  assign {HA_cout_134,HA_out_134}=REGS_372+REGS_373;
  assign {HA_cout_135,HA_out_135}=REGS_374+REGS_375;
  assign {HA_cout_136,HA_out_136}=REGS_376+REGS_377;
  assign {HA_cout_137,HA_out_137}=REGS_378+REGS_379;
  assign {HA_cout_138,HA_out_138}=REGS_380+REGS_381;


  always @(*)
  begin
      REGS_0=inp_0[0];
      REGS_1=HA_out_0;
      REGS_2=HA_out_16;
      REGS_3=HA_cout_16;
      REGS_4=FA_cout_176;
      REGS_5=FA_cout_177;
      REGS_6=FA_cout_178;
      REGS_7=FA_cout_179;
      REGS_8=FA_cout_180;
      REGS_9=FA_cout_181;
      REGS_10=FA_cout_182;
      REGS_11=FA_cout_183;
      REGS_12=FA_cout_184;
      REGS_13=FA_cout_185;
      REGS_14=FA_cout_186;
      REGS_15=FA_cout_187;
      REGS_16=FA_cout_188;
      REGS_17=FA_cout_189;
      REGS_18=FA_cout_190;
      REGS_19=FA_cout_191;
      REGS_20=FA_cout_192;
      REGS_21=FA_cout_193;
      REGS_22=FA_cout_194;
      REGS_23=FA_cout_195;
      REGS_24=FA_cout_196;
      REGS_25=FA_cout_197;
      REGS_26=FA_out_176;
      REGS_27=FA_out_177;
      REGS_28=FA_out_178;
      REGS_29=FA_out_179;
      REGS_30=FA_out_180;
      REGS_31=FA_out_181;
      REGS_32=FA_out_182;
      REGS_33=FA_out_183;
      REGS_34=FA_out_184;
      REGS_35=FA_out_185;
      REGS_36=FA_out_186;
      REGS_37=FA_out_187;
      REGS_38=FA_out_188;
      REGS_39=FA_out_189;
      REGS_40=FA_out_190;
      REGS_41=FA_out_191;
      REGS_42=FA_out_192;
      REGS_43=FA_out_193;
      REGS_44=FA_out_194;
      REGS_45=FA_out_195;
      REGS_46=FA_out_196;
      REGS_47=FA_out_197;
      REGS_48=FA_out_198;
      REGS_49=FA_cout_198;
      REGS_50=FA_out_199;
      REGS_51=FA_cout_199;
      REGS_52=FA_out_200;
      REGS_53=FA_cout_200;
      REGS_54=FA_out_24;
      REGS_55=HA_out_17;
      REGS_56=HA_cout_17;
      REGS_57=HA_cout_18;
      REGS_58=FA_cout_201;
      REGS_59=FA_cout_202;
      REGS_60=FA_cout_203;
      REGS_61=FA_cout_204;
      REGS_62=FA_cout_205;
      REGS_63=FA_cout_206;
      REGS_64=FA_cout_207;
      REGS_65=FA_cout_208;
      REGS_66=FA_cout_209;
      REGS_67=FA_cout_210;
      REGS_68=FA_cout_211;
      REGS_69=FA_cout_212;
      REGS_70=FA_cout_213;
      REGS_71=FA_cout_214;
      REGS_72=FA_cout_215;
      REGS_73=FA_cout_216;
      REGS_74=FA_cout_217;
      REGS_75=FA_out_218;
      REGS_76=FA_cout_218;
      REGS_77=HA_out_18;
      REGS_78=FA_out_201;
      REGS_79=FA_out_202;
      REGS_80=FA_out_203;
      REGS_81=FA_out_204;
      REGS_82=FA_out_205;
      REGS_83=FA_out_206;
      REGS_84=FA_out_207;
      REGS_85=FA_out_208;
      REGS_86=FA_out_209;
      REGS_87=FA_out_210;
      REGS_88=FA_out_211;
      REGS_89=FA_out_212;
      REGS_90=FA_out_213;
      REGS_91=FA_out_214;
      REGS_92=FA_out_215;
      REGS_93=FA_out_216;
      REGS_94=FA_out_217;
      REGS_95=FA_out_219;
      REGS_96=FA_cout_219;
      REGS_97=FA_out_220;
      REGS_98=FA_cout_220;
      REGS_99=FA_out_221;
      REGS_100=FA_cout_221;
      REGS_101=FA_out_222;
      REGS_102=FA_cout_222;
      REGS_103=FA_out_223;
      REGS_104=FA_cout_223;
      REGS_105=FA_out_224;
      REGS_106=FA_cout_224;
      REGS_107=FA_out_225;
      REGS_108=FA_cout_225;
      REGS_109=FA_out_226;
      REGS_110=FA_cout_226;
      REGS_111=inp_9[0];
      REGS_112=HA_out_3;
      REGS_113=HA_out_19;
      REGS_114=HA_cout_19;
      REGS_115=FA_cout_227;
      REGS_116=FA_cout_228;
      REGS_117=FA_cout_229;
      REGS_118=FA_cout_230;
      REGS_119=FA_cout_231;
      REGS_120=FA_cout_232;
      REGS_121=FA_cout_233;
      REGS_122=FA_cout_234;
      REGS_123=FA_cout_235;
      REGS_124=FA_cout_236;
      REGS_125=FA_cout_237;
      REGS_126=FA_cout_238;
      REGS_127=FA_cout_239;
      REGS_128=FA_out_240;
      REGS_129=FA_cout_240;
      REGS_130=FA_out_241;
      REGS_131=FA_cout_241;
      REGS_132=FA_out_227;
      REGS_133=FA_out_228;
      REGS_134=FA_out_229;
      REGS_135=FA_out_230;
      REGS_136=FA_out_231;
      REGS_137=FA_out_232;
      REGS_138=FA_out_233;
      REGS_139=FA_out_234;
      REGS_140=FA_out_235;
      REGS_141=FA_out_236;
      REGS_142=FA_out_237;
      REGS_143=FA_out_238;
      REGS_144=FA_out_239;
      REGS_145=FA_out_242;
      REGS_146=FA_cout_242;
      REGS_147=FA_out_243;
      REGS_148=FA_cout_243;
      REGS_149=FA_out_244;
      REGS_150=FA_cout_244;
      REGS_151=FA_out_245;
      REGS_152=FA_cout_245;
      REGS_153=FA_out_246;
      REGS_154=FA_cout_246;
      REGS_155=FA_out_247;
      REGS_156=FA_cout_247;
      REGS_157=FA_out_248;
      REGS_158=FA_cout_248;
      REGS_159=FA_out_249;
      REGS_160=FA_cout_249;
      REGS_161=FA_out_250;
      REGS_162=FA_cout_250;
      REGS_163=FA_out_96;
      REGS_164=HA_out_20;
      REGS_165=HA_cout_20;
      REGS_166=HA_cout_21;
      REGS_167=FA_cout_251;
      REGS_168=FA_cout_252;
      REGS_169=FA_cout_253;
      REGS_170=FA_cout_254;
      REGS_171=FA_cout_255;
      REGS_172=FA_cout_256;
      REGS_173=FA_cout_257;
      REGS_174=FA_cout_258;
      REGS_175=FA_out_259;
      REGS_176=FA_cout_259;
      REGS_177=FA_out_260;
      REGS_178=FA_cout_260;
      REGS_179=FA_out_261;
      REGS_180=FA_cout_261;
      REGS_181=HA_out_21;
      REGS_182=FA_out_251;
      REGS_183=FA_out_252;
      REGS_184=FA_out_253;
      REGS_185=FA_out_254;
      REGS_186=FA_out_255;
      REGS_187=FA_out_256;
      REGS_188=FA_out_257;
      REGS_189=FA_out_258;
      REGS_190=FA_out_262;
      REGS_191=FA_cout_262;
      REGS_192=FA_out_263;
      REGS_193=FA_cout_263;
      REGS_194=FA_out_264;
      REGS_195=FA_cout_264;
      REGS_196=FA_out_265;
      REGS_197=FA_cout_265;
      REGS_198=FA_out_266;
      REGS_199=FA_cout_266;
      REGS_200=FA_out_267;
      REGS_201=FA_cout_267;
      REGS_202=FA_out_268;
      REGS_203=FA_cout_268;
      REGS_204=FA_out_269;
      REGS_205=FA_cout_269;
      REGS_206=FA_out_270;
      REGS_207=FA_cout_270;
      REGS_208=FA_out_271;
      REGS_209=FA_cout_271;
      REGS_210=FA_out_272;
      REGS_211=FA_cout_272;
      REGS_212=FA_out_273;
      REGS_213=FA_cout_273;
      REGS_214=FA_out_274;
      REGS_215=FA_cout_274;
      REGS_216=FA_out_275;
      REGS_217=FA_cout_275;
      REGS_218=FA_out_276;
      REGS_219=FA_cout_276;
      REGS_220=FA_out_277;
      REGS_221=FA_cout_277;
      REGS_222=inp_18[0];
      REGS_223=HA_out_6;
      REGS_224=HA_out_22;
      REGS_225=HA_cout_22;
      REGS_226=FA_cout_278;
      REGS_227=FA_cout_279;
      REGS_228=FA_cout_280;
      REGS_229=FA_cout_281;
      REGS_230=FA_out_282;
      REGS_231=FA_cout_282;
      REGS_232=FA_out_283;
      REGS_233=FA_cout_283;
      REGS_234=FA_out_284;
      REGS_235=FA_cout_284;
      REGS_236=FA_out_285;
      REGS_237=FA_cout_285;
      REGS_238=FA_out_278;
      REGS_239=FA_out_279;
      REGS_240=FA_out_280;
      REGS_241=FA_out_281;
      REGS_242=FA_out_286;
      REGS_243=FA_cout_286;
      REGS_244=FA_out_287;
      REGS_245=FA_cout_287;
      REGS_246=FA_out_288;
      REGS_247=FA_cout_288;
      REGS_248=FA_out_289;
      REGS_249=FA_cout_289;
      REGS_250=FA_out_290;
      REGS_251=FA_cout_290;
      REGS_252=HA_out_23;
      REGS_253=HA_cout_23;
      REGS_254=FA_out_291;
      REGS_255=FA_cout_291;
      REGS_256=HA_out_24;
      REGS_257=HA_cout_24;
      REGS_258=FA_out_292;
      REGS_259=FA_cout_292;
      REGS_260=HA_out_25;
      REGS_261=HA_cout_25;
      REGS_262=HA_out_26;
      REGS_263=HA_cout_26;
      REGS_264=FA_out_171;
      REGS_265=HA_out_27;
      REGS_266=HA_cout_27;
      REGS_267=FA_out_174;
      REGS_268=HA_out_28;
      REGS_269=HA_cout_28;
      REGS_270=FA_out_168;
      REGS_271=HA_out_8;
      REGS_272=HA_out_29;
      REGS_273=HA_cout_29;
      REGS_274=HA_out_11;
      REGS_275=HA_out_30;
      REGS_276=HA_cout_30;
      REGS_277=HA_out_14;
      REGS_278=HA_out_31;
      REGS_279=HA_cout_31;
      REGS_280=inp_23[2];
      REGS_281=inp_23[11];
      REGS_282=inp_23[20];
      REGS_283=REGS_0;
      REGS_284=REGS_1;
      REGS_285=REGS_2;
      REGS_286=HA_out_32;
      REGS_287=HA_out_49;
      REGS_288=HA_out_65;
      REGS_289=HA_out_83;
      REGS_290=HA_cout_83;
      REGS_291=HA_cout_84;
      REGS_292=HA_cout_85;
      REGS_293=HA_cout_86;
      REGS_294=HA_cout_87;
      REGS_295=HA_cout_88;
      REGS_296=HA_cout_89;
      REGS_297=HA_cout_90;
      REGS_298=HA_cout_91;
      REGS_299=FA_cout_455;
      REGS_300=FA_cout_456;
      REGS_301=FA_cout_457;
      REGS_302=FA_cout_458;
      REGS_303=FA_cout_459;
      REGS_304=FA_cout_460;
      REGS_305=FA_cout_461;
      REGS_306=FA_cout_462;
      REGS_307=FA_cout_463;
      REGS_308=FA_cout_464;
      REGS_309=FA_cout_465;
      REGS_310=FA_cout_466;
      REGS_311=FA_cout_467;
      REGS_312=FA_cout_468;
      REGS_313=HA_out_84;
      REGS_314=HA_out_85;
      REGS_315=HA_out_86;
      REGS_316=HA_out_87;
      REGS_317=HA_out_88;
      REGS_318=HA_out_89;
      REGS_319=HA_out_90;
      REGS_320=HA_out_91;
      REGS_321=FA_out_455;
      REGS_322=FA_out_456;
      REGS_323=FA_out_457;
      REGS_324=FA_out_458;
      REGS_325=FA_out_459;
      REGS_326=FA_out_460;
      REGS_327=FA_out_461;
      REGS_328=FA_out_462;
      REGS_329=FA_out_463;
      REGS_330=FA_out_464;
      REGS_331=FA_out_465;
      REGS_332=FA_out_466;
      REGS_333=FA_out_467;
      REGS_334=FA_out_468;
      REGS_335=FA_out_469;
      REGS_336=FA_cout_469;
      REGS_337=FA_out_470;
      REGS_338=FA_cout_470;
      REGS_339=FA_out_471;
      REGS_340=FA_cout_471;
      REGS_341=FA_out_472;
      REGS_342=FA_cout_472;
      REGS_343=FA_out_473;
      REGS_344=FA_cout_473;
      REGS_345=FA_out_474;
      REGS_346=FA_cout_474;
      REGS_347=FA_out_475;
      REGS_348=FA_cout_475;
      REGS_349=HA_out_71;
      REGS_350=HA_out_72;
      REGS_351=HA_out_73;
      REGS_352=FA_out_446;
      REGS_353=FA_out_447;
      REGS_354=FA_out_448;
      REGS_355=HA_out_74;
      REGS_356=HA_out_92;
      REGS_357=HA_cout_92;
      REGS_358=FA_out_410;
      REGS_359=HA_out_93;
      REGS_360=HA_cout_93;
      REGS_361=HA_out_94;
      REGS_362=HA_cout_94;
      REGS_363=HA_out_95;
      REGS_364=HA_cout_95;
      REGS_365=HA_out_96;
      REGS_366=HA_cout_96;
      REGS_367=HA_out_97;
      REGS_368=HA_cout_97;
      REGS_369=HA_out_98;
      REGS_370=HA_cout_98;
      REGS_371=HA_out_99;
      REGS_372=HA_cout_99;
      REGS_373=HA_out_100;
      REGS_374=HA_cout_100;
      REGS_375=HA_out_101;
      REGS_376=HA_cout_101;
      REGS_377=HA_out_102;
      REGS_378=HA_cout_102;
      REGS_379=HA_out_103;
      REGS_380=HA_cout_103;
      REGS_381=HA_out_104;
      REGS_382=HA_cout_104;
  end


endmodule

