/*
Copyright 2022-2024 Goran Dakov, D.O.B. 11 January 1983, lives in Bristol UK in 2024

Licensed under GPL v3 or commercial license.

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

(* align_width=C,A_out/2,B_out/2 align_height=R *) module icompr(clk,clkEn,R,C,A_out,B_out,and1,is_sig,sig,sm_sig);
  input pwire clk;
  input pwire clkEn;
  input pwire [64:0] R;
  input pwire [64:0] C;
  output pwire [127:0] A_out;
  output pwire [127:0] B_out;
  input pwire and1;
  input pwire sm_sig;
  input pwire sig;
  input pwire is_sig;
  (* register *) reg REGS_0;
  (* register *) reg REGS_1;
  (* register *) reg REGS_2;
  (* register *) reg REGS_3;
  (* register *) reg REGS_4;
  (* register *) reg REGS_5;
  (* register *) reg REGS_6;
  (* register *) reg REGS_7;
  (* register *) reg REGS_8;
  (* register *) reg REGS_9;
  (* register *) reg REGS_10;
  (* register *) reg REGS_11;
  (* register *) reg REGS_12;
  (* register *) reg REGS_13;
  (* register *) reg REGS_14;
  (* register *) reg REGS_15;
  (* register *) reg REGS_16;
  (* register *) reg REGS_17;
  (* register *) reg REGS_18;
  (* register *) reg REGS_19;
  (* register *) reg REGS_20;
  (* register *) reg REGS_21;
  (* register *) reg REGS_22;
  (* register *) reg REGS_23;
  (* register *) reg REGS_24;
  (* register *) reg REGS_25;
  (* register *) reg REGS_26;
  (* register *) reg REGS_27;
  (* register *) reg REGS_28;
  (* register *) reg REGS_29;
  (* register *) reg REGS_30;
  (* register *) reg REGS_31;
  (* register *) reg REGS_32;
  (* register *) reg REGS_33;
  (* register *) reg REGS_34;
  (* register *) reg REGS_35;
  (* register *) reg REGS_36;
  (* register *) reg REGS_37;
  (* register *) reg REGS_38;
  (* register *) reg REGS_39;
  (* register *) reg REGS_40;
  (* register *) reg REGS_41;
  (* register *) reg REGS_42;
  (* register *) reg REGS_43;
  (* register *) reg REGS_44;
  (* register *) reg REGS_45;
  (* register *) reg REGS_46;
  (* register *) reg REGS_47;
  (* register *) reg REGS_48;
  (* register *) reg REGS_49;
  (* register *) reg REGS_50;
  (* register *) reg REGS_51;
  (* register *) reg REGS_52;
  (* register *) reg REGS_53;
  (* register *) reg REGS_54;
  (* register *) reg REGS_55;
  (* register *) reg REGS_56;
  (* register *) reg REGS_57;
  (* register *) reg REGS_58;
  (* register *) reg REGS_59;
  (* register *) reg REGS_60;
  (* register *) reg REGS_61;
  (* register *) reg REGS_62;
  (* register *) reg REGS_63;
  (* register *) reg REGS_64;
  (* register *) reg REGS_65;
  (* register *) reg REGS_66;
  (* register *) reg REGS_67;
  (* register *) reg REGS_68;
  (* register *) reg REGS_69;
  (* register *) reg REGS_70;
  (* register *) reg REGS_71;
  (* register *) reg REGS_72;
  (* register *) reg REGS_73;
  (* register *) reg REGS_74;
  (* register *) reg REGS_75;
  (* register *) reg REGS_76;
  (* register *) reg REGS_77;
  (* register *) reg REGS_78;
  (* register *) reg REGS_79;
  (* register *) reg REGS_80;
  (* register *) reg REGS_81;
  (* register *) reg REGS_82;
  (* register *) reg REGS_83;
  (* register *) reg REGS_84;
  (* register *) reg REGS_85;
  (* register *) reg REGS_86;
  (* register *) reg REGS_87;
  (* register *) reg REGS_88;
  (* register *) reg REGS_89;
  (* register *) reg REGS_90;
  (* register *) reg REGS_91;
  (* register *) reg REGS_92;
  (* register *) reg REGS_93;
  (* register *) reg REGS_94;
  (* register *) reg REGS_95;
  (* register *) reg REGS_96;
  (* register *) reg REGS_97;
  (* register *) reg REGS_98;
  (* register *) reg REGS_99;
  (* register *) reg REGS_100;
  (* register *) reg REGS_101;
  (* register *) reg REGS_102;
  (* register *) reg REGS_103;
  (* register *) reg REGS_104;
  (* register *) reg REGS_105;
  (* register *) reg REGS_106;
  (* register *) reg REGS_107;
  (* register *) reg REGS_108;
  (* register *) reg REGS_109;
  (* register *) reg REGS_110;
  (* register *) reg REGS_111;
  (* register *) reg REGS_112;
  (* register *) reg REGS_113;
  (* register *) reg REGS_114;
  (* register *) reg REGS_115;
  (* register *) reg REGS_116;
  (* register *) reg REGS_117;
  (* register *) reg REGS_118;
  (* register *) reg REGS_119;
  (* register *) reg REGS_120;
  (* register *) reg REGS_121;
  (* register *) reg REGS_122;
  (* register *) reg REGS_123;
  (* register *) reg REGS_124;
  (* register *) reg REGS_125;
  (* register *) reg REGS_126;
  (* register *) reg REGS_127;
  (* register *) reg REGS_128;
  (* register *) reg REGS_129;
  (* register *) reg REGS_130;
  (* register *) reg REGS_131;
  (* register *) reg REGS_132;
  (* register *) reg REGS_133;
  (* register *) reg REGS_134;
  (* register *) reg REGS_135;
  (* register *) reg REGS_136;
  (* register *) reg REGS_137;
  (* register *) reg REGS_138;
  (* register *) reg REGS_139;
  (* register *) reg REGS_140;
  (* register *) reg REGS_141;
  (* register *) reg REGS_142;
  (* register *) reg REGS_143;
  (* register *) reg REGS_144;
  (* register *) reg REGS_145;
  (* register *) reg REGS_146;
  (* register *) reg REGS_147;
  (* register *) reg REGS_148;
  (* register *) reg REGS_149;
  (* register *) reg REGS_150;
  (* register *) reg REGS_151;
  (* register *) reg REGS_152;
  (* register *) reg REGS_153;
  (* register *) reg REGS_154;
  (* register *) reg REGS_155;
  (* register *) reg REGS_156;
  (* register *) reg REGS_157;
  (* register *) reg REGS_158;
  (* register *) reg REGS_159;
  (* register *) reg REGS_160;
  (* register *) reg REGS_161;
  (* register *) reg REGS_162;
  (* register *) reg REGS_163;
  (* register *) reg REGS_164;
  (* register *) reg REGS_165;
  (* register *) reg REGS_166;
  (* register *) reg REGS_167;
  (* register *) reg REGS_168;
  (* register *) reg REGS_169;
  (* register *) reg REGS_170;
  (* register *) reg REGS_171;
  (* register *) reg REGS_172;
  (* register *) reg REGS_173;
  (* register *) reg REGS_174;
  (* register *) reg REGS_175;
  (* register *) reg REGS_176;
  (* register *) reg REGS_177;
  (* register *) reg REGS_178;
  (* register *) reg REGS_179;
  (* register *) reg REGS_180;
  (* register *) reg REGS_181;
  (* register *) reg REGS_182;
  (* register *) reg REGS_183;
  (* register *) reg REGS_184;
  (* register *) reg REGS_185;
  (* register *) reg REGS_186;
  (* register *) reg REGS_187;
  (* register *) reg REGS_188;
  (* register *) reg REGS_189;
  (* register *) reg REGS_190;
  (* register *) reg REGS_191;
  (* register *) reg REGS_192;
  (* register *) reg REGS_193;
  (* register *) reg REGS_194;
  (* register *) reg REGS_195;
  (* register *) reg REGS_196;
  (* register *) reg REGS_197;
  (* register *) reg REGS_198;
  (* register *) reg REGS_199;
  (* register *) reg REGS_200;
  (* register *) reg REGS_201;
  (* register *) reg REGS_202;
  (* register *) reg REGS_203;
  (* register *) reg REGS_204;
  (* register *) reg REGS_205;
  (* register *) reg REGS_206;
  (* register *) reg REGS_207;
  (* register *) reg REGS_208;
  (* register *) reg REGS_209;
  (* register *) reg REGS_210;
  (* register *) reg REGS_211;
  (* register *) reg REGS_212;
  (* register *) reg REGS_213;
  (* register *) reg REGS_214;
  (* register *) reg REGS_215;
  (* register *) reg REGS_216;
  (* register *) reg REGS_217;
  (* register *) reg REGS_218;
  (* register *) reg REGS_219;
  (* register *) reg REGS_220;
  (* register *) reg REGS_221;
  (* register *) reg REGS_222;
  (* register *) reg REGS_223;
  (* register *) reg REGS_224;
  (* register *) reg REGS_225;
  (* register *) reg REGS_226;
  (* register *) reg REGS_227;
  (* register *) reg REGS_228;
  (* register *) reg REGS_229;
  (* register *) reg REGS_230;
  (* register *) reg REGS_231;
  (* register *) reg REGS_232;
  (* register *) reg REGS_233;
  (* register *) reg REGS_234;
  (* register *) reg REGS_235;
  (* register *) reg REGS_236;
  (* register *) reg REGS_237;
  (* register *) reg REGS_238;
  (* register *) reg REGS_239;
  (* register *) reg REGS_240;
  (* register *) reg REGS_241;
  (* register *) reg REGS_242;
  (* register *) reg REGS_243;
  (* register *) reg REGS_244;
  (* register *) reg REGS_245;
  (* register *) reg REGS_246;
  (* register *) reg REGS_247;
  (* register *) reg REGS_248;
  (* register *) reg REGS_249;
  (* register *) reg REGS_250;
  (* register *) reg REGS_251;
  (* register *) reg REGS_252;
  (* register *) reg REGS_253;
  (* register *) reg REGS_254;
  (* register *) reg REGS_255;
  (* register *) reg REGS_256;
  (* register *) reg REGS_257;
  (* register *) reg REGS_258;
  (* register *) reg REGS_259;
  (* register *) reg REGS_260;
  (* register *) reg REGS_261;
  (* register *) reg REGS_262;
  (* register *) reg REGS_263;
  (* register *) reg REGS_264;
  (* register *) reg REGS_265;
  (* register *) reg REGS_266;
  (* register *) reg REGS_267;
  (* register *) reg REGS_268;
  (* register *) reg REGS_269;
  (* register *) reg REGS_270;
  (* register *) reg REGS_271;
  (* register *) reg REGS_272;
  (* register *) reg REGS_273;
  (* register *) reg REGS_274;
  (* register *) reg REGS_275;
  (* register *) reg REGS_276;
  (* register *) reg REGS_277;
  (* register *) reg REGS_278;
  (* register *) reg REGS_279;
  (* register *) reg REGS_280;
  (* register *) reg REGS_281;
  (* register *) reg REGS_282;
  (* register *) reg REGS_283;
  (* register *) reg REGS_284;
  (* register *) reg REGS_285;
  (* register *) reg REGS_286;
  (* register *) reg REGS_287;
  (* register *) reg REGS_288;
  (* register *) reg REGS_289;
  (* register *) reg REGS_290;
  (* register *) reg REGS_291;
  (* register *) reg REGS_292;
  (* register *) reg REGS_293;
  (* register *) reg REGS_294;
  (* register *) reg REGS_295;
  (* register *) reg REGS_296;
  (* register *) reg REGS_297;
  (* register *) reg REGS_298;
  (* register *) reg REGS_299;
  (* register *) reg REGS_300;
  (* register *) reg REGS_301;
  (* register *) reg REGS_302;
  (* register *) reg REGS_303;
  (* register *) reg REGS_304;
  (* register *) reg REGS_305;
  (* register *) reg REGS_306;
  (* register *) reg REGS_307;
  (* register *) reg REGS_308;
  (* register *) reg REGS_309;
  (* register *) reg REGS_310;
  (* register *) reg REGS_311;
  (* register *) reg REGS_312;
  (* register *) reg REGS_313;
  (* register *) reg REGS_314;
  (* register *) reg REGS_315;
  (* register *) reg REGS_316;
  (* register *) reg REGS_317;
  (* register *) reg REGS_318;
  (* register *) reg REGS_319;
  (* register *) reg REGS_320;
  (* register *) reg REGS_321;
  (* register *) reg REGS_322;
  (* register *) reg REGS_323;
  (* register *) reg REGS_324;
  (* register *) reg REGS_325;
  (* register *) reg REGS_326;
  (* register *) reg REGS_327;
  (* register *) reg REGS_328;
  (* register *) reg REGS_329;
  (* register *) reg REGS_330;
  (* register *) reg REGS_331;
  (* register *) reg REGS_332;
  (* register *) reg REGS_333;
  (* register *) reg REGS_334;
  (* register *) reg REGS_335;
  (* register *) reg REGS_336;
  (* register *) reg REGS_337;
  (* register *) reg REGS_338;
  (* register *) reg REGS_339;
  (* register *) reg REGS_340;
  (* register *) reg REGS_341;
  (* register *) reg REGS_342;
  (* register *) reg REGS_343;
  (* register *) reg REGS_344;
  (* register *) reg REGS_345;
  (* register *) reg REGS_346;
  (* register *) reg REGS_347;
  (* register *) reg REGS_348;
  (* register *) reg REGS_349;
  (* register *) reg REGS_350;
  (* register *) reg REGS_351;
  (* register *) reg REGS_352;
  (* register *) reg REGS_353;
  (* register *) reg REGS_354;
  (* register *) reg REGS_355;
  (* register *) reg REGS_356;
  (* register *) reg REGS_357;
  (* register *) reg REGS_358;
  (* register *) reg REGS_359;
  (* register *) reg REGS_360;
  (* register *) reg REGS_361;
  (* register *) reg REGS_362;
  (* register *) reg REGS_363;
  (* register *) reg REGS_364;
  (* register *) reg REGS_365;
  (* register *) reg REGS_366;
  (* register *) reg REGS_367;
  (* register *) reg REGS_368;
  (* register *) reg REGS_369;
  (* register *) reg REGS_370;
  (* register *) reg REGS_371;
  (* register *) reg REGS_372;
  (* register *) reg REGS_373;
  (* register *) reg REGS_374;
  (* register *) reg REGS_375;
  (* register *) reg REGS_376;
  (* register *) reg REGS_377;
  (* register *) reg REGS_378;
  (* register *) reg REGS_379;
  (* register *) reg REGS_380;
  (* register *) reg REGS_381;
  (* register *) reg REGS_382;
  (* register *) reg REGS_383;
  (* register *) reg REGS_384;
  (* register *) reg REGS_385;
  (* register *) reg REGS_386;
  (* register *) reg REGS_387;
  (* register *) reg REGS_388;
  (* register *) reg REGS_389;
  (* register *) reg REGS_390;
  (* register *) reg REGS_391;
  (* register *) reg REGS_392;
  (* register *) reg REGS_393;
  (* register *) reg REGS_394;
  (* register *) reg REGS_395;
  (* register *) reg REGS_396;
  (* register *) reg REGS_397;
  (* register *) reg REGS_398;
  (* register *) reg REGS_399;
  (* register *) reg REGS_400;
  (* register *) reg REGS_401;
  (* register *) reg REGS_402;
  (* register *) reg REGS_403;
  (* register *) reg REGS_404;
  (* register *) reg REGS_405;
  (* register *) reg REGS_406;
  (* register *) reg REGS_407;
  (* register *) reg REGS_408;
  (* register *) reg REGS_409;
  (* register *) reg REGS_410;
  (* register *) reg REGS_411;
  (* register *) reg REGS_412;
  (* register *) reg REGS_413;
  (* register *) reg REGS_414;
  (* register *) reg REGS_415;
  (* register *) reg REGS_416;
  (* register *) reg REGS_417;
  (* register *) reg REGS_418;
  (* register *) reg REGS_419;
  (* register *) reg REGS_420;
  (* register *) reg REGS_421;
  (* register *) reg REGS_422;
  (* register *) reg REGS_423;
  (* register *) reg REGS_424;
  (* register *) reg REGS_425;
  (* register *) reg REGS_426;
  (* register *) reg REGS_427;
  (* register *) reg REGS_428;
  (* register *) reg REGS_429;
  (* register *) reg REGS_430;
  (* register *) reg REGS_431;
  (* register *) reg REGS_432;
  (* register *) reg REGS_433;
  (* register *) reg REGS_434;
  (* register *) reg REGS_435;
  (* register *) reg REGS_436;
  (* register *) reg REGS_437;
  (* register *) reg REGS_438;
  (* register *) reg REGS_439;
  (* register *) reg REGS_440;
  (* register *) reg REGS_441;
  (* register *) reg REGS_442;
  (* register *) reg REGS_443;
  (* register *) reg REGS_444;
  (* register *) reg REGS_445;
  (* register *) reg REGS_446;
  (* register *) reg REGS_447;
  (* register *) reg REGS_448;
  (* register *) reg REGS_449;
  (* register *) reg REGS_450;
  (* register *) reg REGS_451;
  (* register *) reg REGS_452;
  (* register *) reg REGS_453;
  (* register *) reg REGS_454;
  (* register *) reg REGS_455;
  (* register *) reg REGS_456;
  (* register *) reg REGS_457;
  (* register *) reg REGS_458;
  (* register *) reg REGS_459;
  (* register *) reg REGS_460;
  (* register *) reg REGS_461;
  (* register *) reg REGS_462;
  (* register *) reg REGS_463;
  (* register *) reg REGS_464;
  (* register *) reg REGS_465;
  (* register *) reg REGS_466;
  (* register *) reg REGS_467;
  (* register *) reg REGS_468;
  (* register *) reg REGS_469;
  (* register *) reg REGS_470;
  (* register *) reg REGS_471;
  (* register *) reg REGS_472;
  (* register *) reg REGS_473;
  (* register *) reg REGS_474;
  (* register *) reg REGS_475;
  (* register *) reg REGS_476;
  (* register *) reg REGS_477;
  (* register *) reg REGS_478;
  (* register *) reg REGS_479;
  (* register *) reg REGS_480;
  (* register *) reg REGS_481;
  (* register *) reg REGS_482;
  (* register *) reg REGS_483;
  (* register *) reg REGS_484;
  (* register *) reg REGS_485;
  (* register *) reg REGS_486;
  (* register *) reg REGS_487;
  (* register *) reg REGS_488;
  (* register *) reg REGS_489;
  (* register *) reg REGS_490;
  (* register *) reg REGS_491;
  (* register *) reg REGS_492;
  (* register *) reg REGS_493;
  (* register *) reg REGS_494;
  (* register *) reg REGS_495;
  (* register *) reg REGS_496;
  (* register *) reg REGS_497;
  (* register *) reg REGS_498;
  (* register *) reg REGS_499;
  (* register *) reg REGS_500;
  (* register *) reg REGS_501;
  (* register *) reg REGS_502;
  (* register *) reg REGS_503;
  (* register *) reg REGS_504;
  (* register *) reg REGS_505;
  (* register *) reg REGS_506;
  (* register *) reg REGS_507;
  (* register *) reg REGS_508;
  (* register *) reg REGS_509;
  (* register *) reg REGS_510;
  (* register *) reg REGS_511;
  (* register *) reg REGS_512;
  (* register *) reg REGS_513;
  (* register *) reg REGS_514;
  (* register *) reg REGS_515;
  (* register *) reg REGS_516;
  (* register *) reg REGS_517;
  (* register *) reg REGS_518;
  (* register *) reg REGS_519;
  (* register *) reg REGS_520;
  (* register *) reg REGS_521;
  (* register *) reg REGS_522;
  (* register *) reg REGS_523;
  (* register *) reg REGS_524;
  (* register *) reg REGS_525;
  (* register *) reg REGS_526;
  (* register *) reg REGS_527;
  (* register *) reg REGS_528;
  (* register *) reg REGS_529;
  (* register *) reg REGS_530;
  (* register *) reg REGS_531;
  (* register *) reg REGS_532;
  (* register *) reg REGS_533;
  (* register *) reg REGS_534;
  (* register *) reg REGS_535;
  (* register *) reg REGS_536;
  (* register *) reg REGS_537;
  (* register *) reg REGS_538;
  (* register *) reg REGS_539;
  (* register *) reg REGS_540;
  (* register *) reg REGS_541;
  (* register *) reg REGS_542;
  (* register *) reg REGS_543;
  (* register *) reg REGS_544;
  (* register *) reg REGS_545;
  (* register *) reg REGS_546;
  (* register *) reg REGS_547;
  (* register *) reg REGS_548;
  (* register *) reg REGS_549;
  (* register *) reg REGS_550;
  (* register *) reg REGS_551;
  (* register *) reg REGS_552;
  (* register *) reg REGS_553;
  (* register *) reg REGS_554;
  (* register *) reg REGS_555;
  (* register *) reg REGS_556;
  (* register *) reg REGS_557;
  (* register *) reg REGS_558;
  (* register *) reg REGS_559;
  (* register *) reg REGS_560;
  (* register *) reg REGS_561;
  (* register *) reg REGS_562;
  (* register *) reg REGS_563;
  (* register *) reg REGS_564;
  (* register *) reg REGS_565;
  (* register *) reg REGS_566;
  (* register *) reg REGS_567;
  (* register *) reg REGS_568;
  (* register *) reg REGS_569;
  (* register *) reg REGS_570;
  (* register *) reg REGS_571;
  (* register *) reg REGS_572;
  (* register *) reg REGS_573;
  (* register *) reg REGS_574;
  (* register *) reg REGS_575;
  (* register *) reg REGS_576;
  (* register *) reg REGS_577;
  (* register *) reg REGS_578;
  (* register *) reg REGS_579;
  (* register *) reg REGS_580;
  (* register *) reg REGS_581;
  (* register *) reg REGS_582;
  (* register *) reg REGS_583;
  (* register *) reg REGS_584;
  (* register *) reg REGS_585;
  (* register *) reg REGS_586;
  (* register *) reg REGS_587;
  (* register *) reg REGS_588;
  (* register *) reg REGS_589;
  (* register *) reg REGS_590;
  (* register *) reg REGS_591;
  (* register *) reg REGS_592;
  (* register *) reg REGS_593;
  (* register *) reg REGS_594;
  (* register *) reg REGS_595;
  (* register *) reg REGS_596;
  (* register *) reg REGS_597;
  (* register *) reg REGS_598;
  (* register *) reg REGS_599;
  (* register *) reg REGS_600;
  (* register *) reg REGS_601;
  (* register *) reg REGS_602;
  (* register *) reg REGS_603;
  (* register *) reg REGS_604;
  (* register *) reg REGS_605;
  (* register *) reg REGS_606;
  (* register *) reg REGS_607;
  (* register *) reg REGS_608;
  (* register *) reg REGS_609;
  (* register *) reg REGS_610;
  (* register *) reg REGS_611;
  (* register *) reg REGS_612;
  (* register *) reg REGS_613;
  (* register *) reg REGS_614;
  (* register *) reg REGS_615;
  (* register *) reg REGS_616;
  (* register *) reg REGS_617;
  (* register *) reg REGS_618;
  (* register *) reg REGS_619;
  (* register *) reg REGS_620;
  (* register *) reg REGS_621;
  (* register *) reg REGS_622;
  (* register *) reg REGS_623;
  (* register *) reg REGS_624;
  (* register *) reg REGS_625;
  (* register *) reg REGS_626;
  (* register *) reg REGS_627;
  (* register *) reg REGS_628;
  (* register *) reg REGS_629;
  (* register *) reg REGS_630;
  (* register *) reg REGS_631;
  (* register *) reg REGS_632;
  (* register *) reg REGS_633;
  (* register *) reg REGS_634;
  (* register *) reg REGS_635;
  (* register *) reg REGS_636;
  (* register *) reg REGS_637;
  (* register *) reg REGS_638;
  (* register *) reg REGS_639;
  (* register *) reg REGS_640;
  (* register *) reg REGS_641;
  (* register *) reg REGS_642;
  (* register *) reg REGS_643;
  (* register *) reg REGS_644;
  (* register *) reg REGS_645;
  (* register *) reg REGS_646;
  (* register *) reg REGS_647;
  (* register *) reg REGS_648;
  (* register *) reg REGS_649;
  (* register *) reg REGS_650;
  (* register *) reg REGS_651;
  (* register *) reg REGS_652;
  (* register *) reg REGS_653;
  (* register *) reg REGS_654;
  (* register *) reg REGS_655;
  (* register *) reg REGS_656;
  (* register *) reg REGS_657;
  (* register *) reg REGS_658;
  (* register *) reg REGS_659;
  (* register *) reg REGS_660;
  (* register *) reg REGS_661;
  (* register *) reg REGS_662;
  (* register *) reg REGS_663;
  (* register *) reg REGS_664;
  (* register *) reg REGS_665;
  (* register *) reg REGS_666;
  (* register *) reg REGS_667;
  (* register *) reg REGS_668;
  (* register *) reg REGS_669;
  (* register *) reg REGS_670;
  (* register *) reg REGS_671;
  (* register *) reg REGS_672;
  (* register *) reg REGS_673;
  (* register *) reg REGS_674;
  (* register *) reg REGS_675;
  (* register *) reg REGS_676;
  (* register *) reg REGS_677;
  (* register *) reg REGS_678;
  (* register *) reg REGS_679;
  (* register *) reg REGS_680;
  (* register *) reg REGS_681;
  (* register *) reg REGS_682;
  (* register *) reg REGS_683;
  (* register *) reg REGS_684;
  (* register *) reg REGS_685;
  (* register *) reg REGS_686;
  (* register *) reg REGS_687;
  (* register *) reg REGS_688;
  (* register *) reg REGS_689;
  (* register *) reg REGS_690;
  (* register *) reg REGS_691;
  (* register *) reg REGS_692;
  (* register *) reg REGS_693;
  (* register *) reg REGS_694;
  (* register *) reg REGS_695;
  (* register *) reg REGS_696;
  (* register *) reg REGS_697;
  (* register *) reg REGS_698;
  (* register *) reg REGS_699;
  (* register *) reg REGS_700;
  (* register *) reg REGS_701;
  (* register *) reg REGS_702;
  (* register *) reg REGS_703;
  (* register *) reg REGS_704;
  (* register *) reg REGS_705;
  (* register *) reg REGS_706;
  (* register *) reg REGS_707;
  (* register *) reg REGS_708;
  (* register *) reg REGS_709;
  (* register *) reg REGS_710;
  (* register *) reg REGS_711;
  (* register *) reg REGS_712;
  (* register *) reg REGS_713;
  (* register *) reg REGS_714;
  (* register *) reg REGS_715;
  (* register *) reg REGS_716;
  (* register *) reg REGS_717;
  (* register *) reg REGS_718;
  (* register *) reg REGS_719;
  (* register *) reg REGS_720;
  (* register *) reg REGS_721;
  (* register *) reg REGS_722;
  (* register *) reg REGS_723;
  (* register *) reg REGS_724;
  (* register *) reg REGS_725;
  (* register *) reg REGS_726;
  (* register *) reg REGS_727;
  (* register *) reg REGS_728;
  (* register *) reg REGS_729;
  (* register *) reg REGS_730;
  (* register *) reg REGS_731;
  (* register *) reg REGS_732;
  (* register *) reg REGS_733;
  (* register *) reg REGS_734;
  (* register *) reg REGS_735;
  (* register *) reg REGS_736;
  (* register *) reg REGS_737;
  (* register *) reg REGS_738;
  (* register *) reg REGS_739;
  (* register *) reg REGS_740;
  (* register *) reg REGS_741;
  (* register *) reg REGS_742;
  (* register *) reg REGS_743;
  (* register *) reg REGS_744;
  (* register *) reg REGS_745;
  (* register *) reg REGS_746;
  (* register *) reg REGS_747;
  (* register *) reg REGS_748;
  (* register *) reg REGS_749;
  (* register *) reg REGS_750;
  (* register *) reg REGS_751;
  (* register *) reg REGS_752;
  (* register *) reg REGS_753;
  (* register *) reg REGS_754;
  (* register *) reg REGS_755;
  (* register *) reg REGS_756;
  (* register *) reg REGS_757;
  (* register *) reg REGS_758;
  (* register *) reg REGS_759;
  (* register *) reg REGS_760;
  (* register *) reg REGS_761;
  (* register *) reg REGS_762;
  (* register *) reg REGS_763;
  (* register *) reg REGS_764;
  (* register *) reg REGS_765;
  (* register *) reg REGS_766;
  (* register *) reg REGS_767;
  (* register *) reg REGS_768;
  (* register *) reg REGS_769;
  (* register *) reg REGS_770;
  (* register *) reg REGS_771;
  (* register *) reg REGS_772;
  (* register *) reg REGS_773;
  (* register *) reg REGS_774;
  (* register *) reg REGS_775;
  (* register *) reg REGS_776;
  (* register *) reg REGS_777;
  (* register *) reg REGS_778;
  (* register *) reg REGS_779;
  (* register *) reg REGS_780;
  (* register *) reg REGS_781;
  (* register *) reg REGS_782;
  (* register *) reg REGS_783;
  (* register *) reg REGS_784;
  (* register *) reg REGS_785;
  (* register *) reg REGS_786;
  (* register *) reg REGS_787;
  (* register *) reg REGS_788;
  (* register *) reg REGS_789;
  (* register *) reg REGS_790;
  (* register *) reg REGS_791;
  (* register *) reg REGS_792;
  (* register *) reg REGS_793;
  (* register *) reg REGS_794;
  (* register *) reg REGS_795;
  (* register *) reg REGS_796;
  (* register *) reg REGS_797;
  (* register *) reg REGS_798;
  (* register *) reg REGS_799;
  (* register *) reg REGS_800;
  (* register *) reg REGS_801;
  (* register *) reg REGS_802;
  (* register *) reg REGS_803;
  (* register *) reg REGS_804;
  (* register *) reg REGS_805;
  (* register *) reg REGS_806;
  (* register *) reg REGS_807;
  (* register *) reg REGS_808;
  (* register *) reg REGS_809;
  (* register *) reg REGS_810;
  (* register *) reg REGS_811;
  (* register *) reg REGS_812;
  (* register *) reg REGS_813;
  (* register *) reg REGS_814;
  (* register *) reg REGS_815;
  (* register *) reg REGS_816;
  (* register *) reg REGS_817;
  (* register *) reg REGS_818;
  (* register *) reg REGS_819;
  (* register *) reg REGS_820;
  (* register *) reg REGS_821;
  (* register *) reg REGS_822;
  (* register *) reg REGS_823;
  (* register *) reg REGS_824;
  (* register *) reg REGS_825;
  (* register *) reg REGS_826;
  (* register *) reg REGS_827;
  (* register *) reg REGS_828;
  (* register *) reg REGS_829;
  (* register *) reg REGS_830;
  (* register *) reg REGS_831;
  (* register *) reg REGS_832;
  (* register *) reg REGS_833;
  (* register *) reg REGS_834;
  (* register *) reg REGS_835;
  (* register *) reg REGS_836;
  (* register *) reg REGS_837;
  (* register *) reg REGS_838;
  (* register *) reg REGS_839;
  (* register *) reg REGS_840;
  (* register *) reg REGS_841;
  (* register *) reg REGS_842;
  (* register *) reg REGS_843;
  (* register *) reg REGS_844;
  (* register *) reg REGS_845;
  (* register *) reg REGS_846;
  (* register *) reg REGS_847;
  (* register *) reg REGS_848;
  (* register *) reg REGS_849;
  (* register *) reg REGS_850;
  (* register *) reg REGS_851;
  (* register *) reg REGS_852;
  (* register *) reg REGS_853;
  (* register *) reg REGS_854;
  (* register *) reg REGS_855;
  (* register *) reg REGS_856;
  (* register *) reg REGS_857;
  (* register *) reg REGS_858;
  (* register *) reg REGS_859;
  (* register *) reg REGS_860;
  (* register *) reg REGS_861;
  (* register *) reg REGS_862;
  (* register *) reg REGS_863;
  (* register *) reg REGS_864;
  (* register *) reg REGS_865;
  (* register *) reg REGS_866;
  (* register *) reg REGS_867;
  (* register *) reg REGS_868;
  (* register *) reg REGS_869;
  (* register *) reg REGS_870;
  (* register *) reg REGS_871;
  (* register *) reg REGS_872;
  (* register *) reg REGS_873;
  (* register *) reg REGS_874;
  (* register *) reg REGS_875;
  (* register *) reg REGS_876;
  (* register *) reg REGS_877;
  (* register *) reg REGS_878;
  (* register *) reg REGS_879;
  (* register *) reg REGS_880;
  (* register *) reg REGS_881;
  (* register *) reg REGS_882;
  (* register *) reg REGS_883;
  (* register *) reg REGS_884;
  (* register *) reg REGS_885;
  (* register *) reg REGS_886;
  (* register *) reg REGS_887;
  (* register *) reg REGS_888;
  (* register *) reg REGS_889;
  (* register *) reg REGS_890;
  (* register *) reg REGS_891;
  (* register *) reg REGS_892;
  (* register *) reg REGS_893;
  (* register *) reg REGS_894;
  (* register *) reg REGS_895;
  (* register *) reg REGS_896;
  (* register *) reg REGS_897;
  (* register *) reg REGS_898;
  (* register *) reg REGS_899;
  (* register *) reg REGS_900;
  (* register *) reg REGS_901;
  (* register *) reg REGS_902;
  (* register *) reg REGS_903;
  (* register *) reg REGS_904;
  (* register *) reg REGS_905;
  (* register *) reg REGS_906;
  (* register *) reg REGS_907;
  (* register *) reg REGS_908;
  (* register *) reg REGS_909;
  (* register *) reg REGS_910;
  (* register *) reg REGS_911;
  (* register *) reg REGS_912;
  (* register *) reg REGS_913;
  (* register *) reg REGS_914;
  (* register *) reg REGS_915;
  (* register *) reg REGS_916;
  (* register *) reg REGS_917;
  (* register *) reg REGS_918;
  (* register *) reg REGS_919;
  (* register *) reg REGS_920;
  (* register *) reg REGS_921;
  (* register *) reg REGS_922;
  (* register *) reg REGS_923;
  (* register *) reg REGS_924;
  (* register *) reg REGS_925;
  (* register *) reg REGS_926;
  (* register *) reg REGS_927;
  (* register *) reg REGS_928;
  (* register *) reg REGS_929;
  (* register *) reg REGS_930;
  (* register *) reg REGS_931;
  (* register *) reg REGS_932;
  (* register *) reg REGS_933;
  (* register *) reg REGS_934;
  (* register *) reg REGS_935;
  (* register *) reg REGS_936;
  (* register *) reg REGS_937;
  (* register *) reg REGS_938;
  (* register *) reg REGS_939;
  (* register *) reg REGS_940;
  (* register *) reg REGS_941;
  (* register *) reg REGS_942;
  (* register *) reg REGS_943;
  (* register *) reg REGS_944;
  (* register *) reg REGS_945;
  (* register *) reg REGS_946;
  (* register *) reg REGS_947;
  (* register *) reg REGS_948;
  (* register *) reg REGS_949;
  (* register *) reg REGS_950;
  (* register *) reg REGS_951;
  (* register *) reg REGS_952;
  (* register *) reg REGS_953;
  (* register *) reg REGS_954;
  (* register *) reg REGS_955;
  (* register *) reg REGS_956;
  (* register *) reg REGS_957;
  (* register *) reg REGS_958;
  (* register *) reg REGS_959;
  (* register *) reg REGS_960;
  (* register *) reg REGS_961;
  (* register *) reg REGS_962;
  (* register *) reg REGS_963;
  (* register *) reg REGS_964;
  (* register *) reg REGS_965;
  (* register *) reg REGS_966;
  (* register *) reg REGS_967;
  (* register *) reg REGS_968;
  (* register *) reg REGS_969;
  (* register *) reg REGS_970;
  (* register *) reg REGS_971;
  (* register *) reg REGS_972;
  (* register *) reg REGS_973;
  (* register *) reg REGS_974;
  (* register *) reg REGS_975;
  (* register *) reg REGS_976;
  (* register *) reg REGS_977;
  (* register *) reg REGS_978;
  (* register *) reg REGS_979;
  (* register *) reg REGS_980;
  (* register *) reg REGS_981;
  (* register *) reg REGS_982;
  (* register *) reg REGS_983;
  (* register *) reg REGS_984;
  (* register *) reg REGS_985;
  (* register *) reg REGS_986;
  (* register *) reg REGS_987;
  (* register *) reg REGS_988;
  (* register *) reg REGS_989;
  (* register *) reg REGS_990;
  (* register *) reg REGS_991;
  (* register *) reg REGS_992;
  (* register *) reg REGS_993;
  (* register *) reg REGS_994;
  (* register *) reg REGS_995;
  (* register *) reg REGS_996;
  (* register *) reg REGS_997;
  (* register *) reg REGS_998;
  (* register *) reg REGS_999;
  (* register *) reg REGS_1000;
  (* register *) reg REGS_1001;
  (* register *) reg REGS_1002;
  (* register *) reg REGS_1003;
  (* register *) reg REGS_1004;
  (* register *) reg REGS_1005;
  (* register *) reg REGS_1006;
  (* register *) reg REGS_1007;
  (* register *) reg REGS_1008;
  (* register *) reg REGS_1009;
  (* register *) reg REGS_1010;
  (* register *) reg REGS_1011;
  (* register *) reg REGS_1012;
  (* register *) reg REGS_1013;
  (* register *) reg REGS_1014;
  (* register *) reg REGS_1015;
  (* register *) reg REGS_1016;
  (* register *) reg REGS_1017;
  (* register *) reg REGS_1018;
  (* register *) reg REGS_1019;
  (* register *) reg REGS_1020;
  (* register *) reg REGS_1021;
  (* register *) reg REGS_1022;
  (* register *) reg REGS_1023;
  (* register *) reg REGS_1024;
  (* register *) reg REGS_1025;
  (* register *) reg REGS_1026;
  (* register *) reg REGS_1027;
  (* register *) reg REGS_1028;
  (* register *) reg REGS_1029;
  (* register *) reg REGS_1030;
  (* register *) reg REGS_1031;
  (* register *) reg REGS_1032;
  (* register *) reg REGS_1033;
  (* register *) reg REGS_1034;
  (* register *) reg REGS_1035;
  (* register *) reg REGS_1036;
  (* register *) reg REGS_1037;
  (* register *) reg REGS_1038;
  (* register *) reg REGS_1039;
  (* register *) reg REGS_1040;
  (* register *) reg REGS_1041;
  (* register *) reg REGS_1042;
  (* register *) reg REGS_1043;
  (* register *) reg REGS_1044;
  (* register *) reg REGS_1045;
  (* register *) reg REGS_1046;
  (* register *) reg REGS_1047;
  (* register *) reg REGS_1048;
  (* register *) reg REGS_1049;
  (* register *) reg REGS_1050;
  (* register *) reg REGS_1051;
  (* register *) reg REGS_1052;
  (* register *) reg REGS_1053;
  (* register *) reg REGS_1054;
  (* register *) reg REGS_1055;
  (* register *) reg REGS_1056;
  (* register *) reg REGS_1057;
  (* register *) reg REGS_1058;
  (* register *) reg REGS_1059;
  (* register *) reg REGS_1060;
  (* register *) reg REGS_1061;
  (* register *) reg REGS_1062;
  (* register *) reg REGS_1063;
  (* register *) reg REGS_1064;
  (* register *) reg REGS_1065;
  (* register *) reg REGS_1066;
  (* register *) reg REGS_1067;
  (* register *) reg REGS_1068;
  (* register *) reg REGS_1069;
  (* register *) reg REGS_1070;
  (* register *) reg REGS_1071;
  (* register *) reg REGS_1072;
  (* register *) reg REGS_1073;
  (* register *) reg REGS_1074;
  (* register *) reg REGS_1075;
  (* register *) reg REGS_1076;
  (* register *) reg REGS_1077;
  (* register *) reg REGS_1078;
  (* register *) reg REGS_1079;
  (* register *) reg REGS_1080;
  (* register *) reg REGS_1081;
  (* register *) reg REGS_1082;
  (* register *) reg REGS_1083;
  (* register *) reg REGS_1084;
  (* register *) reg REGS_1085;
  (* register *) reg REGS_1086;
  (* register *) reg REGS_1087;
  (* register *) reg REGS_1088;
  (* register *) reg REGS_1089;
  (* register *) reg REGS_1090;
  (* register *) reg REGS_1091;
  (* register *) reg REGS_1092;
  (* register *) reg REGS_1093;
  (* register *) reg REGS_1094;
  (* register *) reg REGS_1095;
  (* register *) reg REGS_1096;
  (* register *) reg REGS_1097;
  (* register *) reg REGS_1098;
  (* register *) reg REGS_1099;
  (* register *) reg REGS_1100;
  (* register *) reg REGS_1101;
  (* register *) reg REGS_1102;
  (* register *) reg REGS_1103;
  (* register *) reg REGS_1104;
  (* register *) reg REGS_1105;
  (* register *) reg REGS_1106;
  (* register *) reg REGS_1107;
  (* register *) reg REGS_1108;
  (* register *) reg REGS_1109;
  (* register *) reg REGS_1110;
  (* register *) reg REGS_1111;
  (* register *) reg REGS_1112;
  (* register *) reg REGS_1113;
  (* register *) reg REGS_1114;
  (* register *) reg REGS_1115;
  (* register *) reg REGS_1116;
  (* register *) reg REGS_1117;
  (* register *) reg REGS_1118;
  (* register *) reg REGS_1119;
  (* register *) reg REGS_1120;
  (* register *) reg REGS_1121;
  (* register *) reg REGS_1122;
  (* register *) reg REGS_1123;
  (* register *) reg REGS_1124;
  (* register *) reg REGS_1125;
  (* register *) reg REGS_1126;
  (* register *) reg REGS_1127;
  (* register *) reg REGS_1128;
  (* register *) reg REGS_1129;
  (* register *) reg REGS_1130;
  (* register *) reg REGS_1131;
  (* register *) reg REGS_1132;
  (* register *) reg REGS_1133;
  (* register *) reg REGS_1134;
  (* register *) reg REGS_1135;
  (* register *) reg REGS_1136;
  (* register *) reg REGS_1137;
  (* register *) reg REGS_1138;
  (* register *) reg REGS_1139;
  (* register *) reg REGS_1140;
  (* register *) reg REGS_1141;
  (* register *) reg REGS_1142;
  (* register *) reg REGS_1143;
  (* register *) reg REGS_1144;
  (* register *) reg REGS_1145;
  (* register *) reg REGS_1146;
  (* register *) reg REGS_1147;
  (* register *) reg REGS_1148;
  (* register *) reg REGS_1149;
  (* register *) reg REGS_1150;
  (* register *) reg REGS_1151;
  (* register *) reg REGS_1152;
  (* register *) reg REGS_1153;
  (* register *) reg REGS_1154;
  (* register *) reg REGS_1155;
  (* register *) reg REGS_1156;
  (* register *) reg REGS_1157;
  (* register *) reg REGS_1158;
  (* register *) reg REGS_1159;
  (* register *) reg REGS_1160;
  (* register *) reg REGS_1161;
  (* register *) reg REGS_1162;
  (* register *) reg REGS_1163;
  (* register *) reg REGS_1164;
  (* register *) reg REGS_1165;
  (* register *) reg REGS_1166;
  (* register *) reg REGS_1167;
  (* register *) reg REGS_1168;
  (* register *) reg REGS_1169;
  (* register *) reg REGS_1170;
  (* register *) reg REGS_1171;
  (* register *) reg REGS_1172;
  (* register *) reg REGS_1173;
  (* register *) reg REGS_1174;
  (* register *) reg REGS_1175;
  (* register *) reg REGS_1176;
  (* register *) reg REGS_1177;
  (* register *) reg REGS_1178;
  (* register *) reg REGS_1179;
  (* register *) reg REGS_1180;
  (* register *) reg REGS_1181;
  (* register *) reg REGS_1182;
  (* register *) reg REGS_1183;
  (* register *) reg REGS_1184;
  (* register *) reg REGS_1185;
  (* register *) reg REGS_1186;
  (* register *) reg REGS_1187;
  (* register *) reg REGS_1188;
  (* register *) reg REGS_1189;
  (* register *) reg REGS_1190;
  (* register *) reg REGS_1191;
  (* register *) reg REGS_1192;
  (* register *) reg REGS_1193;
  (* register *) reg REGS_1194;
  (* register *) reg REGS_1195;
  (* register *) reg REGS_1196;
  (* register *) reg REGS_1197;
  (* register *) reg REGS_1198;
  (* register *) reg REGS_1199;
  (* register *) reg REGS_1200;
  (* register *) reg REGS_1201;
  (* register *) reg REGS_1202;
  (* register *) reg REGS_1203;
  (* register *) reg REGS_1204;
  (* register *) reg REGS_1205;
  (* register *) reg REGS_1206;
  (* register *) reg REGS_1207;
  (* register *) reg REGS_1208;
  (* register *) reg REGS_1209;
  (* register *) reg REGS_1210;
  (* register *) reg REGS_1211;
  (* register *) reg REGS_1212;
  (* register *) reg REGS_1213;
  (* register *) reg REGS_1214;
  (* register *) reg REGS_1215;
  (* register *) reg REGS_1216;
  (* register *) reg REGS_1217;
  (* register *) reg REGS_1218;
  (* register *) reg REGS_1219;
  (* register *) reg REGS_1220;
  (* register *) reg REGS_1221;
  (* register *) reg REGS_1222;
  (* register *) reg REGS_1223;
  (* register *) reg REGS_1224;
  (* register *) reg REGS_1225;
  (* register *) reg REGS_1226;
  (* register *) reg REGS_1227;
  (* register *) reg REGS_1228;
  (* register *) reg REGS_1229;
  (* register *) reg REGS_1230;
  (* register *) reg REGS_1231;
  (* register *) reg REGS_1232;
  (* register *) reg REGS_1233;
  (* register *) reg REGS_1234;
  (* register *) reg REGS_1235;
  (* register *) reg REGS_1236;
  (* register *) reg REGS_1237;
  (* register *) reg REGS_1238;
  (* register *) reg REGS_1239;
  (* register *) reg REGS_1240;
  (* register *) reg REGS_1241;
  (* register *) reg REGS_1242;
  (* register *) reg REGS_1243;
  (* register *) reg REGS_1244;
  (* register *) reg REGS_1245;
  (* register *) reg REGS_1246;
  (* register *) reg REGS_1247;
  (* register *) reg REGS_1248;
  (* register *) reg REGS_1249;
  (* register *) reg REGS_1250;
  (* register *) reg REGS_1251;
  (* register *) reg REGS_1252;
  (* register *) reg REGS_1253;
  (* register *) reg REGS_1254;
  (* register *) reg REGS_1255;
  (* register *) reg REGS_1256;
  (* register *) reg REGS_1257;
  (* register *) reg REGS_1258;
  (* register *) reg REGS_1259;
  (* register *) reg REGS_1260;
  (* register *) reg REGS_1261;
  (* register *) reg REGS_1262;
  (* register *) reg REGS_1263;
  (* register *) reg REGS_1264;
  (* register *) reg REGS_1265;
  (* register *) reg REGS_1266;
  (* register *) reg REGS_1267;
  (* register *) reg REGS_1268;
  (* register *) reg REGS_1269;
  (* register *) reg REGS_1270;
  (* register *) reg REGS_1271;
  (* register *) reg REGS_1272;
  (* register *) reg REGS_1273;
  (* register *) reg REGS_1274;
  (* register *) reg REGS_1275;
  (* register *) reg REGS_1276;
  (* register *) reg REGS_1277;
  (* register *) reg REGS_1278;
  (* register *) reg REGS_1279;
  (* register *) reg REGS_1280;
  (* register *) reg REGS_1281;
  (* register *) reg REGS_1282;
  (* register *) reg REGS_1283;
  (* register *) reg REGS_1284;
  (* register *) reg REGS_1285;
  (* register *) reg REGS_1286;
  (* register *) reg REGS_1287;
  (* register *) reg REGS_1288;
  (* register *) reg REGS_1289;
  (* register *) reg REGS_1290;
  (* register *) reg REGS_1291;
  (* register *) reg REGS_1292;
  (* register *) reg REGS_1293;
  (* register *) reg REGS_1294;
  (* register *) reg REGS_1295;
  (* register *) reg REGS_1296;
  (* register *) reg REGS_1297;
  (* register *) reg REGS_1298;
  (* register *) reg REGS_1299;
  (* register *) reg REGS_1300;
  (* register *) reg REGS_1301;
  (* register *) reg REGS_1302;
  (* register *) reg REGS_1303;
  (* register *) reg REGS_1304;
  (* register *) reg REGS_1305;
  (* register *) reg REGS_1306;
  (* register *) reg REGS_1307;
  (* register *) reg REGS_1308;
  (* register *) reg REGS_1309;
  (* register *) reg REGS_1310;
  (* register *) reg REGS_1311;
  (* register *) reg REGS_1312;
  (* register *) reg REGS_1313;
  (* register *) reg REGS_1314;
  (* register *) reg REGS_1315;
  (* register *) reg REGS_1316;
  (* register *) reg REGS_1317;
  (* register *) reg REGS_1318;
  (* register *) reg REGS_1319;
  (* register *) reg REGS_1320;
  (* register *) reg REGS_1321;
  (* register *) reg REGS_1322;
  (* register *) reg REGS_1323;
  (* register *) reg REGS_1324;
  (* register *) reg REGS_1325;
  (* register *) reg REGS_1326;
  (* register *) reg REGS_1327;
  (* register *) reg REGS_1328;
  (* register *) reg REGS_1329;
  (* register *) reg REGS_1330;
  (* register *) reg REGS_1331;
  (* register *) reg REGS_1332;
  (* register *) reg REGS_1333;
  (* register *) reg REGS_1334;
  (* register *) reg REGS_1335;
  (* register *) reg REGS_1336;
  (* register *) reg REGS_1337;
  (* register *) reg REGS_1338;
  (* register *) reg REGS_1339;
  (* register *) reg REGS_1340;
  (* register *) reg REGS_1341;
  (* register *) reg REGS_1342;
  (* register *) reg REGS_1343;
  (* register *) reg REGS_1344;
  (* register *) reg REGS_1345;
  (* register *) reg REGS_1346;
  (* register *) reg REGS_1347;
  (* register *) reg REGS_1348;
  (* register *) reg REGS_1349;
  (* register *) reg REGS_1350;
  (* register *) reg REGS_1351;
  (* register *) reg REGS_1352;
  (* register *) reg REGS_1353;
  (* register *) reg REGS_1354;
  (* register *) reg REGS_1355;
  (* register *) reg REGS_1356;
  (* register *) reg REGS_1357;
  (* register *) reg REGS_1358;
  (* register *) reg REGS_1359;
  (* register *) reg REGS_1360;
  (* register *) reg REGS_1361;
  (* register *) reg REGS_1362;
  (* register *) reg REGS_1363;
  (* register *) reg REGS_1364;
  (* register *) reg REGS_1365;
  (* register *) reg REGS_1366;
  (* register *) reg REGS_1367;
  (* register *) reg REGS_1368;
  (* register *) reg REGS_1369;
  (* register *) reg REGS_1370;
  (* register *) reg REGS_1371;
  (* register *) reg REGS_1372;
  (* register *) reg REGS_1373;
  (* register *) reg REGS_1374;
  (* register *) reg REGS_1375;
  (* register *) reg REGS_1376;
  (* register *) reg REGS_1377;
  (* register *) reg REGS_1378;
  (* register *) reg REGS_1379;
  (* register *) reg REGS_1380;
  (* register *) reg REGS_1381;
  (* register *) reg REGS_1382;
  (* register *) reg REGS_1383;
  (* register *) reg REGS_1384;
  (* register *) reg REGS_1385;
  (* register *) reg REGS_1386;
  (* register *) reg REGS_1387;
  (* register *) reg REGS_1388;
  (* register *) reg REGS_1389;
  (* register *) reg REGS_1390;
  (* register *) reg REGS_1391;
  (* register *) reg REGS_1392;
  (* register *) reg REGS_1393;
  (* register *) reg REGS_1394;
  (* register *) reg REGS_1395;
  (* register *) reg REGS_1396;
  (* register *) reg REGS_1397;
  (* register *) reg REGS_1398;
  (* register *) reg REGS_1399;
  (* register *) reg REGS_1400;
  (* register *) reg REGS_1401;
  (* register *) reg REGS_1402;
  (* register *) reg REGS_1403;
  (* register *) reg REGS_1404;
  (* register *) reg REGS_1405;
  (* register *) reg REGS_1406;
  (* register *) reg REGS_1407;
  (* register *) reg REGS_1408;
  (* register *) reg REGS_1409;
  (* register *) reg REGS_1410;
  (* register *) reg REGS_1411;
  (* register *) reg REGS_1412;
  (* register *) reg REGS_1413;
  (* register *) reg REGS_1414;
  (* register *) reg REGS_1415;
  (* register *) reg REGS_1416;
  (* register *) reg REGS_1417;
  (* register *) reg REGS_1418;
  (* register *) reg REGS_1419;
  (* register *) reg REGS_1420;
  (* register *) reg REGS_1421;
  (* register *) reg REGS_1422;
  (* register *) reg REGS_1423;
  (* register *) reg REGS_1424;
  (* register *) reg REGS_1425;
  (* register *) reg REGS_1426;
  (* register *) reg REGS_1427;
  (* register *) reg REGS_1428;
  (* register *) reg REGS_1429;
  (* register *) reg REGS_1430;
  (* register *) reg REGS_1431;
  (* register *) reg REGS_1432;
  (* register *) reg REGS_1433;
  (* register *) reg REGS_1434;
  (* register *) reg REGS_1435;
  (* register *) reg REGS_1436;
  (* register *) reg REGS_1437;
  (* register *) reg REGS_1438;
  (* register *) reg REGS_1439;
  (* register *) reg REGS_1440;
  (* register *) reg REGS_1441;
  (* register *) reg REGS_1442;
  (* register *) reg REGS_1443;
  (* register *) reg REGS_1444;
  (* register *) reg REGS_1445;
  (* register *) reg REGS_1446;
  (* register *) reg REGS_1447;
  (* register *) reg REGS_1448;
  (* register *) reg REGS_1449;
  (* register *) reg REGS_1450;
  (* register *) reg REGS_1451;
  (* register *) reg REGS_1452;
  (* register *) reg REGS_1453;
  (* register *) reg REGS_1454;
  (* register *) reg REGS_1455;
  (* register *) reg REGS_1456;
  (* register *) reg REGS_1457;
  (* register *) reg REGS_1458;
  (* register *) reg REGS_1459;
  (* register *) reg REGS_1460;
  (* register *) reg REGS_1461;
  (* register *) reg REGS_1462;
  (* register *) reg REGS_1463;
  (* register *) reg REGS_1464;
  (* register *) reg REGS_1465;
  (* register *) reg REGS_1466;
  (* register *) reg REGS_1467;
  (* register *) reg REGS_1468;
  (* register *) reg REGS_1469;
  (* register *) reg REGS_1470;
  (* register *) reg REGS_1471;
  (* register *) reg REGS_1472;
  (* register *) reg REGS_1473;
  (* register *) reg REGS_1474;
  (* register *) reg REGS_1475;
  (* register *) reg REGS_1476;
  (* register *) reg REGS_1477;
  (* register *) reg REGS_1478;
  (* register *) reg REGS_1479;
  (* register *) reg REGS_1480;
  (* register *) reg REGS_1481;
  (* register *) reg REGS_1482;
  (* register *) reg REGS_1483;
  (* register *) reg REGS_1484;
  (* register *) reg REGS_1485;
  (* register *) reg REGS_1486;
  (* register *) reg REGS_1487;
  (* register *) reg REGS_1488;
  (* register *) reg REGS_1489;
  (* register *) reg REGS_1490;
  (* register *) reg REGS_1491;
  (* register *) reg REGS_1492;
  (* register *) reg REGS_1493;
  (* register *) reg REGS_1494;
  (* register *) reg REGS_1495;
  (* register *) reg REGS_1496;
  (* register *) reg REGS_1497;
  (* register *) reg REGS_1498;
  (* register *) reg REGS_1499;
  (* register *) reg REGS_1500;
  (* register *) reg REGS_1501;
  (* register *) reg REGS_1502;
  (* register *) reg REGS_1503;
  (* register *) reg REGS_1504;
  (* register *) reg REGS_1505;
  (* register *) reg REGS_1506;
  (* register *) reg REGS_1507;
  (* register *) reg REGS_1508;
  (* register *) reg REGS_1509;
  (* register *) reg REGS_1510;
  (* register *) reg REGS_1511;
  (* register *) reg REGS_1512;
  (* register *) reg REGS_1513;
  (* register *) reg REGS_1514;
  (* register *) reg REGS_1515;
  (* register *) reg REGS_1516;
  (* register *) reg REGS_1517;
  (* register *) reg REGS_1518;
  (* register *) reg REGS_1519;
  (* register *) reg REGS_1520;
  (* register *) reg REGS_1521;
  (* register *) reg REGS_1522;
  (* register *) reg REGS_1523;
  (* register *) reg REGS_1524;
  (* register *) reg REGS_1525;
  (* register *) reg REGS_1526;
  (* register *) reg REGS_1527;
  (* register *) reg REGS_1528;
  (* register *) reg REGS_1529;
  (* register *) reg REGS_1530;
  (* register *) reg REGS_1531;
  (* register *) reg REGS_1532;
  (* register *) reg REGS_1533;
  (* register *) reg REGS_1534;
  (* register *) reg REGS_1535;
  (* register *) reg REGS_1536;
  (* register *) reg REGS_1537;
  (* register *) reg REGS_1538;
  (* register *) reg REGS_1539;
  (* register *) reg REGS_1540;
  (* register *) reg REGS_1541;
  (* register *) reg REGS_1542;
  (* register *) reg REGS_1543;
  (* register *) reg REGS_1544;
  (* register *) reg REGS_1545;
  (* register *) reg REGS_1546;
  (* register *) reg REGS_1547;
  (* register *) reg REGS_1548;
  (* register *) reg REGS_1549;
  (* register *) reg REGS_1550;
  (* register *) reg REGS_1551;
  (* register *) reg REGS_1552;
  (* register *) reg REGS_1553;
  (* register *) reg REGS_1554;
  (* register *) reg REGS_1555;
  (* register *) reg REGS_1556;
  (* register *) reg REGS_1557;
  (* register *) reg REGS_1558;
  (* register *) reg REGS_1559;
  (* register *) reg REGS_1560;
  (* register *) reg REGS_1561;
  (* register *) reg REGS_1562;
  (* register *) reg REGS_1563;
  (* register *) reg REGS_1564;
  (* register *) reg REGS_1565;
  (* register *) reg REGS_1566;
  (* register *) reg REGS_1567;
  (* register *) reg REGS_1568;
  (* register *) reg REGS_1569;
  (* register *) reg REGS_1570;
  (* register *) reg REGS_1571;
  (* register *) reg REGS_1572;
  (* register *) reg REGS_1573;
  (* register *) reg REGS_1574;
  (* register *) reg REGS_1575;
  (* register *) reg REGS_1576;
  (* register *) reg REGS_1577;
  (* register *) reg REGS_1578;
  (* register *) reg REGS_1579;
  (* register *) reg REGS_1580;
  (* register *) reg REGS_1581;
  (* register *) reg REGS_1582;
  (* register *) reg REGS_1583;
  (* register *) reg REGS_1584;
  (* register *) reg REGS_1585;
  (* register *) reg REGS_1586;
  (* register *) reg REGS_1587;
  (* register *) reg REGS_1588;
  (* register *) reg REGS_1589;
  (* register *) reg REGS_1590;
  (* register *) reg REGS_1591;
  (* register *) reg REGS_1592;
  (* register *) reg REGS_1593;
  (* register *) reg REGS_1594;
  (* register *) reg REGS_1595;
  (* register *) reg REGS_1596;
  (* register *) reg REGS_1597;
  (* register *) reg REGS_1598;
  (* register *) reg REGS_1599;
  (* register *) reg REGS_1600;
  (* register *) reg REGS_1601;
  (* register *) reg REGS_1602;
  (* register *) reg REGS_1603;
  (* register *) reg REGS_1604;
  (* register *) reg REGS_1605;
  (* register *) reg REGS_1606;
  (* register *) reg REGS_1607;
  (* register *) reg REGS_1608;
  (* register *) reg REGS_1609;
  (* register *) reg REGS_1610;
  (* register *) reg REGS_1611;
  (* register *) reg REGS_1612;
  (* register *) reg REGS_1613;
  (* register *) reg REGS_1614;
  (* register *) reg REGS_1615;
  (* register *) reg REGS_1616;
  (* register *) reg REGS_1617;
  (* register *) reg REGS_1618;
  (* register *) reg REGS_1619;
  (* register *) reg REGS_1620;
  (* register *) reg REGS_1621;
  (* register *) reg REGS_1622;
  (* register *) reg REGS_1623;
  (* register *) reg REGS_1624;
  (* register *) reg REGS_1625;
  (* register *) reg REGS_1626;
  (* register *) reg REGS_1627;
  (* register *) reg REGS_1628;
  (* register *) reg REGS_1629;
  (* register *) reg REGS_1630;
  (* register *) reg REGS_1631;
  (* register *) reg REGS_1632;
  (* register *) reg REGS_1633;
  (* register *) reg REGS_1634;
  (* register *) reg REGS_1635;
  (* register *) reg REGS_1636;
  (* register *) reg REGS_1637;
  (* register *) reg REGS_1638;
  (* register *) reg REGS_1639;
  (* register *) reg REGS_1640;
  (* register *) reg REGS_1641;
  (* register *) reg REGS_1642;
  (* register *) reg REGS_1643;
  (* register *) reg REGS_1644;
  (* register *) reg REGS_1645;
  (* register *) reg REGS_1646;
  (* register *) reg REGS_1647;
  (* register *) reg REGS_1648;
  (* register *) reg REGS_1649;
  (* register *) reg REGS_1650;
  (* register *) reg REGS_1651;
  (* register *) reg REGS_1652;
  (* register *) reg REGS_1653;
  (* register *) reg REGS_1654;
  (* register *) reg REGS_1655;
  (* register *) reg REGS_1656;
  (* register *) reg REGS_1657;
  (* register *) reg REGS_1658;
  (* register *) reg REGS_1659;
  (* register *) reg REGS_1660;
  (* register *) reg REGS_1661;
  (* register *) reg REGS_1662;
  (* register *) reg REGS_1663;
  (* register *) reg REGS_1664;
  (* register *) reg REGS_1665;
  (* register *) reg REGS_1666;
  (* register *) reg REGS_1667;
  (* register *) reg REGS_1668;
  (* register *) reg REGS_1669;
  (* register *) reg REGS_1670;
  (* register *) reg REGS_1671;
  (* register *) reg REGS_1672;
  (* register *) reg REGS_1673;
  (* register *) reg REGS_1674;
  (* register *) reg REGS_1675;
  (* register *) reg REGS_1676;
  (* register *) reg REGS_1677;
  (* register *) reg REGS_1678;
  (* register *) reg REGS_1679;
  (* register *) reg REGS_1680;
  (* register *) reg REGS_1681;
  (* register *) reg REGS_1682;
  (* register *) reg REGS_1683;
  (* register *) reg REGS_1684;
  (* register *) reg REGS_1685;
  (* register *) reg REGS_1686;
  (* register *) reg REGS_1687;
  (* register *) reg REGS_1688;
  (* register *) reg REGS_1689;
  (* register *) reg REGS_1690;
  (* register *) reg REGS_1691;
  (* register *) reg REGS_1692;
  (* register *) reg REGS_1693;
  (* register *) reg REGS_1694;
  (* register *) reg REGS_1695;
  (* register *) reg REGS_1696;
  (* register *) reg REGS_1697;
  (* register *) reg REGS_1698;
  (* register *) reg REGS_1699;
  (* register *) reg REGS_1700;
  (* register *) reg REGS_1701;
  (* register *) reg REGS_1702;
  (* register *) reg REGS_1703;
  (* register *) reg REGS_1704;
  (* register *) reg REGS_1705;
  (* register *) reg REGS_1706;
  (* register *) reg REGS_1707;
  (* register *) reg REGS_1708;
  (* register *) reg REGS_1709;
  (* register *) reg REGS_1710;
  (* register *) reg REGS_1711;
  (* register *) reg REGS_1712;
  (* register *) reg REGS_1713;
  (* register *) reg REGS_1714;
  (* register *) reg REGS_1715;
  (* register *) reg REGS_1716;
  (* register *) reg REGS_1717;
  (* register *) reg REGS_1718;
  (* register *) reg REGS_1719;
  (* register *) reg REGS_1720;
  (* register *) reg REGS_1721;
  (* register *) reg REGS_1722;
  (* register *) reg REGS_1723;
  (* register *) reg REGS_1724;
  (* register *) reg REGS_1725;
  (* register *) reg REGS_1726;
  (* register *) reg REGS_1727;
  (* register *) reg REGS_1728;
  (* register *) reg REGS_1729;
  (* register *) reg REGS_1730;
  (* register *) reg REGS_1731;
  (* register *) reg REGS_1732;
  (* register *) reg REGS_1733;
  (* register *) reg REGS_1734;
  (* register *) reg REGS_1735;
  (* register *) reg REGS_1736;
  (* register *) reg REGS_1737;
  (* register *) reg REGS_1738;
  (* register *) reg REGS_1739;
  (* register *) reg REGS_1740;
  (* register *) reg REGS_1741;
  (* register *) reg REGS_1742;
  (* register *) reg REGS_1743;
  (* register *) reg REGS_1744;
  (* register *) reg REGS_1745;
  (* register *) reg REGS_1746;
  (* register *) reg REGS_1747;
  (* register *) reg REGS_1748;
  (* register *) reg REGS_1749;
  (* register *) reg REGS_1750;
  (* register *) reg REGS_1751;
  (* register *) reg REGS_1752;
  (* register *) reg REGS_1753;
  (* register *) reg REGS_1754;
  (* register *) reg REGS_1755;
  (* register *) reg REGS_1756;
  (* register *) reg REGS_1757;
  (* register *) reg REGS_1758;
  (* register *) reg REGS_1759;
  (* register *) reg REGS_1760;
  (* register *) reg REGS_1761;
  (* register *) reg REGS_1762;
  (* register *) reg REGS_1763;
  (* register *) reg REGS_1764;
  (* register *) reg REGS_1765;
  (* register *) reg REGS_1766;
  (* register *) reg REGS_1767;
  (* register *) reg REGS_1768;
  (* register *) reg REGS_1769;
  (* register *) reg REGS_1770;
  (* register *) reg REGS_1771;
  (* register *) reg REGS_1772;
  (* register *) reg REGS_1773;
  (* register *) reg REGS_1774;
  (* register *) reg REGS_1775;
  (* register *) reg REGS_1776;
  (* register *) reg REGS_1777;
  (* register *) reg REGS_1778;
  (* register *) reg REGS_1779;
  (* register *) reg REGS_1780;
  (* register *) reg REGS_1781;
  (* register *) reg REGS_1782;
  (* register *) reg REGS_1783;
  (* register *) reg REGS_1784;
  (* register *) reg REGS_1785;
  (* register *) reg REGS_1786;
  (* register *) reg REGS_1787;
  (* register *) reg REGS_1788;
  (* register *) reg REGS_1789;
  (* register *) reg REGS_1790;
  (* register *) reg REGS_1791;
  (* register *) reg REGS_1792;
  (* register *) reg REGS_1793;
  (* register *) reg REGS_1794;
  (* register *) reg REGS_1795;
  (* register *) reg REGS_1796;
  (* register *) reg REGS_1797;
  (* register *) reg REGS_1798;
  (* register *) reg REGS_1799;
  (* register *) reg REGS_1800;
  (* register *) reg REGS_1801;
  (* register *) reg REGS_1802;
  (* register *) reg REGS_1803;
  (* register *) reg REGS_1804;
  (* register *) reg REGS_1805;
  (* register *) reg REGS_1806;
  (* register *) reg REGS_1807;
  (* register *) reg REGS_1808;
  (* register *) reg REGS_1809;
  (* register *) reg REGS_1810;
  (* register *) reg REGS_1811;
  (* register *) reg REGS_1812;
  (* register *) reg REGS_1813;
  (* register *) reg REGS_1814;
  (* register *) reg REGS_1815;
  (* register *) reg REGS_1816;
  (* register *) reg REGS_1817;
  (* register *) reg REGS_1818;
  (* register *) reg REGS_1819;
  (* register *) reg REGS_1820;
  (* register *) reg REGS_1821;
  (* register *) reg REGS_1822;
  (* register *) reg REGS_1823;
  (* register *) reg REGS_1824;
  (* register *) reg REGS_1825;
  (* register *) reg REGS_1826;
  (* register *) reg REGS_1827;
  (* register *) reg REGS_1828;
  (* register *) reg REGS_1829;
  (* register *) reg REGS_1830;
  (* register *) reg REGS_1831;
  (* register *) reg REGS_1832;
  (* register *) reg REGS_1833;
  (* register *) reg REGS_1834;
  (* register *) reg REGS_1835;
  (* register *) reg REGS_1836;
  (* register *) reg REGS_1837;
  (* register *) reg REGS_1838;
  (* register *) reg REGS_1839;
  (* register *) reg REGS_1840;
  (* register *) reg REGS_1841;
  (* register *) reg REGS_1842;
  (* register *) reg REGS_1843;
  (* register *) reg REGS_1844;
  (* register *) reg REGS_1845;
  (* register *) reg REGS_1846;
  (* register *) reg REGS_1847;
  (* register *) reg REGS_1848;
  (* register *) reg REGS_1849;
  (* register *) reg REGS_1850;
  (* register *) reg REGS_1851;
  (* register *) reg REGS_1852;
  (* register *) reg REGS_1853;
  (* register *) reg REGS_1854;
  (* register *) reg REGS_1855;
  (* register *) reg REGS_1856;
  (* register *) reg REGS_1857;
  (* register *) reg REGS_1858;
  (* register *) reg REGS_1859;
  (* register *) reg REGS_1860;
  (* register *) reg REGS_1861;
  (* register *) reg REGS_1862;
  (* register *) reg REGS_1863;
  (* register *) reg REGS_1864;
  (* register *) reg REGS_1865;
  (* register *) reg REGS_1866;
  (* register *) reg REGS_1867;
  (* register *) reg REGS_1868;
  (* register *) reg REGS_1869;
  (* register *) reg REGS_1870;
  (* register *) reg REGS_1871;
  (* register *) reg REGS_1872;
  (* register *) reg REGS_1873;
  (* register *) reg REGS_1874;
  (* register *) reg REGS_1875;
  (* register *) reg REGS_1876;
  (* register *) reg REGS_1877;
  (* register *) reg REGS_1878;
  (* register *) reg REGS_1879;
  (* register *) reg REGS_1880;
  (* register *) reg REGS_1881;
  (* register *) reg REGS_1882;
  (* register *) reg REGS_1883;
  (* register *) reg REGS_1884;
  (* register *) reg REGS_1885;
  (* register *) reg REGS_1886;
  (* register *) reg REGS_1887;
  (* register *) reg REGS_1888;
  (* register *) reg REGS_1889;
  (* register *) reg REGS_1890;
  (* register *) reg REGS_1891;
  (* register *) reg REGS_1892;
  (* register *) reg REGS_1893;
  (* register *) reg REGS_1894;
  (* register *) reg REGS_1895;
  (* register *) reg REGS_1896;
  (* register *) reg REGS_1897;
  (* register *) reg REGS_1898;
  (* register *) reg REGS_1899;
  (* register *) reg REGS_1900;
  (* register *) reg REGS_1901;
  (* register *) reg REGS_1902;
  (* register *) reg REGS_1903;
  (* register *) reg REGS_1904;
  (* register *) reg REGS_1905;
  (* register *) reg REGS_1906;
  (* register *) reg REGS_1907;
  (* register *) reg REGS_1908;
  (* register *) reg REGS_1909;
  (* register *) reg REGS_1910;
  (* register *) reg REGS_1911;
  (* register *) reg REGS_1912;
  (* register *) reg REGS_1913;
  (* register *) reg REGS_1914;
  (* register *) reg REGS_1915;
  (* register *) reg REGS_1916;
  (* register *) reg REGS_1917;
  (* register *) reg REGS_1918;
  (* register *) reg REGS_1919;
  (* register *) reg REGS_1920;
  (* register *) reg REGS_1921;
  (* register *) reg REGS_1922;
  (* register *) reg REGS_1923;
  (* register *) reg REGS_1924;
  (* register *) reg REGS_1925;
  (* register *) reg REGS_1926;
  (* register *) reg REGS_1927;
  (* register *) reg REGS_1928;
  (* register *) reg REGS_1929;
  (* register *) reg REGS_1930;
  (* register *) reg REGS_1931;
  (* register *) reg REGS_1932;
  (* register *) reg REGS_1933;
  (* register *) reg REGS_1934;
  (* register *) reg REGS_1935;
  (* register *) reg REGS_1936;
  (* register *) reg REGS_1937;
  (* register *) reg REGS_1938;
  (* register *) reg REGS_1939;
  (* register *) reg REGS_1940;
  (* register *) reg REGS_1941;
  (* register *) reg REGS_1942;
  (* register *) reg REGS_1943;
  (* register *) reg REGS_1944;
  (* register *) reg REGS_1945;
  (* register *) reg REGS_1946;
  (* register *) reg REGS_1947;
  (* register *) reg REGS_1948;
  (* register *) reg REGS_1949;
  (* register *) reg REGS_1950;
  (* register *) reg REGS_1951;
  (* register *) reg REGS_1952;
  (* register *) reg REGS_1953;
  (* register *) reg REGS_1954;
  (* register *) reg REGS_1955;
  (* register *) reg REGS_1956;
  (* register *) reg REGS_1957;
  (* register *) reg REGS_1958;
  (* register *) reg REGS_1959;
  (* register *) reg REGS_1960;
  (* register *) reg REGS_1961;
  (* register *) reg REGS_1962;
  (* register *) reg REGS_1963;
  (* register *) reg REGS_1964;
  (* register *) reg REGS_1965;
  (* register *) reg REGS_1966;
  (* register *) reg REGS_1967;
  (* register *) reg REGS_1968;
  (* register *) reg REGS_1969;
  (* register *) reg REGS_1970;
  (* register *) reg REGS_1971;
  (* register *) reg REGS_1972;
  (* register *) reg REGS_1973;
  (* register *) reg REGS_1974;
  (* register *) reg REGS_1975;
  (* register *) reg REGS_1976;
  (* register *) reg REGS_1977;
  (* register *) reg REGS_1978;
  (* register *) reg REGS_1979;
  (* register *) reg REGS_1980;
  (* register *) reg REGS_1981;
  (* register *) reg REGS_1982;
  (* register *) reg REGS_1983;
  (* register *) reg REGS_1984;
  (* register *) reg REGS_1985;
  (* register *) reg REGS_1986;
  (* register *) reg REGS_1987;
  (* register *) reg REGS_1988;
  (* register *) reg REGS_1989;
  (* register *) reg REGS_1990;
  (* register *) reg REGS_1991;
  (* register *) reg REGS_1992;
  (* register *) reg REGS_1993;
  (* register *) reg REGS_1994;
  (* register *) reg REGS_1995;
  (* register *) reg REGS_1996;
  (* register *) reg REGS_1997;
  (* register *) reg REGS_1998;
  (* register *) reg REGS_1999;
  (* register *) reg REGS_2000;
  (* register *) reg REGS_2001;
  (* register *) reg REGS_2002;
  (* register *) reg REGS_2003;
  (* register *) reg REGS_2004;
  (* register *) reg REGS_2005;
  (* register *) reg REGS_2006;
  (* register *) reg REGS_2007;
  (* register *) reg REGS_2008;
  (* register *) reg REGS_2009;
  (* register *) reg REGS_2010;
  (* register *) reg REGS_2011;
  (* register *) reg REGS_2012;
  (* register *) reg REGS_2013;
  (* register *) reg REGS_2014;
  (* register *) reg REGS_2015;
  (* register *) reg REGS_2016;
  (* register *) reg REGS_2017;
  (* register *) reg REGS_2018;
  (* register *) reg REGS_2019;
  (* register *) reg REGS_2020;
  (* register *) reg REGS_2021;
  (* register *) reg REGS_2022;
  (* register *) reg REGS_2023;
  (* register *) reg REGS_2024;
  (* register *) reg REGS_2025;
  (* register *) reg REGS_2026;
  (* register *) reg REGS_2027;
  (* register *) reg REGS_2028;
  (* register *) reg REGS_2029;
  (* register *) reg REGS_2030;
  (* register *) reg REGS_2031;
  (* register *) reg REGS_2032;
  (* register *) reg REGS_2033;
  (* register *) reg REGS_2034;
  (* register *) reg REGS_2035;
  (* register *) reg REGS_2036;
  (* register *) reg REGS_2037;
  (* register *) reg REGS_2038;
  (* register *) reg REGS_2039;
  (* register *) reg REGS_2040;
  (* register *) reg REGS_2041;
  (* register *) reg REGS_2042;
  (* register *) reg REGS_2043;
  (* register *) reg REGS_2044;
  (* register *) reg REGS_2045;
  (* register *) reg REGS_2046;
  (* register *) reg REGS_2047;
  (* register *) reg REGS_2048;
  (* register *) reg REGS_2049;
  (* register *) reg REGS_2050;
  (* register *) reg REGS_2051;
  (* register *) reg REGS_2052;
  (* register *) reg REGS_2053;
  (* register *) reg REGS_2054;
  (* register *) reg REGS_2055;
  (* register *) reg REGS_2056;
  (* register *) reg REGS_2057;
  (* register *) reg REGS_2058;
  (* register *) reg REGS_2059;
  (* register *) reg REGS_2060;
  (* register *) reg REGS_2061;
  (* register *) reg REGS_2062;
  (* register *) reg REGS_2063;
  (* register *) reg REGS_2064;
  (* register *) reg REGS_2065;
  (* register *) reg REGS_2066;
  (* register *) reg REGS_2067;
  (* register *) reg REGS_2068;
  (* register *) reg REGS_2069;
  (* register *) reg REGS_2070;
  (* register *) reg REGS_2071;
  (* register *) reg REGS_2072;
  (* register *) reg REGS_2073;
  (* register *) reg REGS_2074;
  (* register *) reg REGS_2075;
  (* register *) reg REGS_2076;
  (* register *) reg REGS_2077;
  (* register *) reg REGS_2078;
  (* register *) reg REGS_2079;
  (* register *) reg REGS_2080;
  (* register *) reg REGS_2081;
  (* register *) reg REGS_2082;
  (* register *) reg REGS_2083;
  (* register *) reg REGS_2084;
  (* register *) reg REGS_2085;
  (* register *) reg REGS_2086;
  (* register *) reg REGS_2087;
  (* register *) reg REGS_2088;
  (* register *) reg REGS_2089;
  (* register *) reg REGS_2090;
  (* register *) reg REGS_2091;
  (* register *) reg REGS_2092;
  (* register *) reg REGS_2093;
  (* register *) reg REGS_2094;
  (* register *) reg REGS_2095;
  (* register *) reg REGS_2096;
  (* register *) reg REGS_2097;
  (* register *) reg REGS_2098;
  (* register *) reg REGS_2099;
  (* register *) reg REGS_2100;
  (* register *) reg REGS_2101;
  (* register *) reg REGS_2102;
  (* register *) reg REGS_2103;
  (* register *) reg REGS_2104;
  (* register *) reg REGS_2105;
  (* register *) reg REGS_2106;
  (* register *) reg REGS_2107;
  (* register *) reg REGS_2108;
  (* register *) reg REGS_2109;
  (* register *) reg REGS_2110;
  (* register *) reg REGS_2111;
  (* register *) reg REGS_2112;
  (* register *) reg REGS_2113;
  (* register *) reg REGS_2114;
  (* register *) reg REGS_2115;
  (* register *) reg REGS_2116;
  (* register *) reg REGS_2117;
  (* register *) reg REGS_2118;
  (* register *) reg REGS_2119;
  (* register *) reg REGS_2120;
  (* register *) reg REGS_2121;
  (* register *) reg REGS_2122;
  (* register *) reg REGS_2123;
  (* register *) reg REGS_2124;
  (* register *) reg REGS_2125;
  (* register *) reg REGS_2126;
  (* register *) reg REGS_2127;
  (* register *) reg REGS_2128;
  (* register *) reg REGS_2129;
  (* register *) reg REGS_2130;
  (* register *) reg REGS_2131;
  (* register *) reg REGS_2132;
  (* register *) reg REGS_2133;
  (* register *) reg REGS_2134;
  (* register *) reg REGS_2135;
  (* register *) reg REGS_2136;
  (* register *) reg REGS_2137;
  (* register *) reg REGS_2138;
  (* register *) reg REGS_2139;
  (* register *) reg REGS_2140;
  (* register *) reg REGS_2141;
  (* register *) reg REGS_2142;
  (* register *) reg REGS_2143;
  (* register *) reg REGS_2144;
  (* register *) reg REGS_2145;
  (* register *) reg REGS_2146;
  (* register *) reg REGS_2147;
  (* register *) reg REGS_2148;
  (* register *) reg REGS_2149;
  (* register *) reg REGS_2150;
  (* register *) reg REGS_2151;
  (* register *) reg REGS_2152;
  (* register *) reg REGS_2153;
  (* register *) reg REGS_2154;
  (* register *) reg REGS_2155;
  (* register *) reg REGS_2156;
  (* register *) reg REGS_2157;
  (* register *) reg REGS_2158;
  (* register *) reg REGS_2159;
  (* register *) reg REGS_2160;
  (* register *) reg REGS_2161;
  (* register *) reg REGS_2162;
  (* register *) reg REGS_2163;
  (* register *) reg REGS_2164;
  (* register *) reg REGS_2165;
  (* register *) reg REGS_2166;
  (* register *) reg REGS_2167;
  (* register *) reg REGS_2168;
  (* register *) reg REGS_2169;
  (* register *) reg REGS_2170;
  (* register *) reg REGS_2171;
  (* register *) reg REGS_2172;
  (* register *) reg REGS_2173;
  (* register *) reg REGS_2174;
  (* register *) reg REGS_2175;
  (* register *) reg REGS_2176;
  (* register *) reg REGS_2177;
  (* register *) reg REGS_2178;
  (* register *) reg REGS_2179;
  (* register *) reg REGS_2180;
  (* register *) reg REGS_2181;
  (* register *) reg REGS_2182;
  (* register *) reg REGS_2183;
  (* register *) reg REGS_2184;
  (* register *) reg REGS_2185;
  (* register *) reg REGS_2186;
  (* register *) reg REGS_2187;
  (* register *) reg REGS_2188;
  (* register *) reg REGS_2189;
  (* register *) reg REGS_2190;
  (* register *) reg REGS_2191;
  (* register *) reg REGS_2192;
  (* register *) reg REGS_2193;
  (* register *) reg REGS_2194;
  (* register *) reg REGS_2195;
  (* register *) reg REGS_2196;
  (* register *) reg REGS_2197;
  (* register *) reg REGS_2198;
  (* register *) reg REGS_2199;
  (* register *) reg REGS_2200;
  (* register *) reg REGS_2201;
  (* register *) reg REGS_2202;
  (* register *) reg REGS_2203;
  (* register *) reg REGS_2204;
  (* register *) reg REGS_2205;
  (* register *) reg REGS_2206;
  (* register *) reg REGS_2207;
  (* register *) reg REGS_2208;
  (* register *) reg REGS_2209;
  (* register *) reg REGS_2210;
  (* register *) reg REGS_2211;
  (* register *) reg REGS_2212;
  (* register *) reg REGS_2213;
  (* register *) reg REGS_2214;
  (* register *) reg REGS_2215;
  (* register *) reg REGS_2216;
  (* register *) reg REGS_2217;
  (* register *) reg REGS_2218;
  (* register *) reg REGS_2219;
  (* register *) reg REGS_2220;
  (* register *) reg REGS_2221;
  (* register *) reg REGS_2222;
  (* register *) reg REGS_2223;
  (* register *) reg REGS_2224;
  (* register *) reg REGS_2225;
  (* register *) reg REGS_2226;
  (* register *) reg REGS_2227;
  (* register *) reg REGS_2228;
  (* register *) reg REGS_2229;
  (* register *) reg REGS_2230;
  (* register *) reg REGS_2231;
  (* register *) reg REGS_2232;
  (* register *) reg REGS_2233;
  (* register *) reg REGS_2234;
  (* register *) reg REGS_2235;
  (* register *) reg REGS_2236;
  (* register *) reg REGS_2237;
  (* register *) reg REGS_2238;
  (* register *) reg REGS_2239;
  (* register *) reg REGS_2240;
  (* register *) reg REGS_2241;
  (* register *) reg REGS_2242;
  (* register *) reg REGS_2243;
  (* register *) reg REGS_2244;
  (* register *) reg REGS_2245;
  (* register *) reg REGS_2246;
  (* register *) reg REGS_2247;
  (* register *) reg REGS_2248;
  (* register *) reg REGS_2249;
  (* register *) reg REGS_2250;
  (* register *) reg REGS_2251;
  (* register *) reg REGS_2252;
  (* register *) reg REGS_2253;
  (* register *) reg REGS_2254;
  (* register *) reg REGS_2255;
  (* register *) reg REGS_2256;
  (* register *) reg REGS_2257;
  (* register *) reg REGS_2258;
  (* register *) reg REGS_2259;
  (* register *) reg REGS_2260;
  (* register *) reg REGS_2261;
  (* register *) reg REGS_2262;
  (* register *) reg REGS_2263;
  (* register *) reg REGS_2264;
  (* register *) reg REGS_2265;
  (* register *) reg REGS_2266;
  (* register *) reg REGS_2267;
  (* register *) reg REGS_2268;
  (* register *) reg REGS_2269;
  (* register *) reg REGS_2270;
  (* register *) reg REGS_2271;
  (* register *) reg REGS_2272;
  (* register *) reg REGS_2273;
  (* register *) reg REGS_2274;
  (* register *) reg REGS_2275;
  (* register *) reg REGS_2276;
  (* register *) reg REGS_2277;
  (* register *) reg REGS_2278;
  (* register *) reg REGS_2279;
  (* register *) reg REGS_2280;
  (* register *) reg REGS_2281;
  (* register *) reg REGS_2282;
  (* register *) reg REGS_2283;
  (* register *) reg REGS_2284;
  (* register *) reg REGS_2285;
  (* register *) reg REGS_2286;
  (* register *) reg REGS_2287;
  (* register *) reg REGS_2288;
  (* register *) reg REGS_2289;
  (* register *) reg REGS_2290;
  (* register *) reg REGS_2291;
  (* register *) reg REGS_2292;
  (* register *) reg REGS_2293;
  (* register *) reg REGS_2294;
  (* register *) reg REGS_2295;
  (* register *) reg REGS_2296;
  (* register *) reg REGS_2297;
  (* register *) reg REGS_2298;
  (* register *) reg REGS_2299;
  (* register *) reg REGS_2300;
  (* register *) reg REGS_2301;
  (* register *) reg REGS_2302;
  (* register *) reg REGS_2303;
  (* register *) reg REGS_2304;
  (* register *) reg REGS_2305;
  (* register *) reg REGS_2306;
  (* register *) reg REGS_2307;
  (* register *) reg REGS_2308;
  (* register *) reg REGS_2309;
  (* register *) reg REGS_2310;
  (* register *) reg REGS_2311;
  (* register *) reg REGS_2312;
  (* register *) reg REGS_2313;
  (* register *) reg REGS_2314;
  (* register *) reg REGS_2315;
  (* register *) reg REGS_2316;
  (* register *) reg REGS_2317;
  (* register *) reg REGS_2318;
  (* register *) reg REGS_2319;
  (* register *) reg REGS_2320;
  (* register *) reg REGS_2321;
  (* register *) reg REGS_2322;
  (* register *) reg REGS_2323;
  (* register *) reg REGS_2324;
  (* register *) reg REGS_2325;
  (* register *) reg REGS_2326;
  (* register *) reg REGS_2327;
  (* register *) reg REGS_2328;
  (* register *) reg REGS_2329;
  (* register *) reg REGS_2330;
  (* register *) reg REGS_2331;
  (* register *) reg REGS_2332;
  (* register *) reg REGS_2333;
  (* register *) reg REGS_2334;
  (* register *) reg REGS_2335;
  (* register *) reg REGS_2336;
  (* register *) reg REGS_2337;
  (* register *) reg REGS_2338;
  (* register *) reg REGS_2339;
  (* register *) reg REGS_2340;
  (* register *) reg REGS_2341;
  (* register *) reg REGS_2342;
  (* register *) reg REGS_2343;
  (* register *) reg REGS_2344;
  (* register *) reg REGS_2345;
  (* register *) reg REGS_2346;
  (* register *) reg REGS_2347;
  (* register *) reg REGS_2348;
  (* register *) reg REGS_2349;
  (* register *) reg REGS_2350;
  (* register *) reg REGS_2351;
  (* register *) reg REGS_2352;
  (* register *) reg REGS_2353;
  (* register *) reg REGS_2354;
  (* register *) reg REGS_2355;
  (* register *) reg REGS_2356;
  (* register *) reg REGS_2357;
  (* register *) reg REGS_2358;
  (* register *) reg REGS_2359;
  (* register *) reg REGS_2360;
  (* register *) reg REGS_2361;
  (* register *) reg REGS_2362;
  (* register *) reg REGS_2363;
  (* register *) reg REGS_2364;
  (* register *) reg REGS_2365;
  (* register *) reg REGS_2366;
  (* register *) reg REGS_2367;
  (* register *) reg REGS_2368;
  (* register *) reg REGS_2369;
  (* register *) reg REGS_2370;
  (* register *) reg REGS_2371;
  (* register *) reg REGS_2372;
  (* register *) reg REGS_2373;
  (* register *) reg REGS_2374;
  (* register *) reg REGS_2375;
  (* register *) reg REGS_2376;
  (* register *) pwire FA_out_0;
  (* register *) pwire FA_out_1;
  (* register *) pwire FA_out_2;
  (* register *) pwire FA_out_3;
  (* register *) pwire FA_out_4;
  (* register *) pwire FA_out_5;
  (* register *) pwire FA_out_6;
  (* register *) pwire FA_out_7;
  (* register *) pwire FA_out_8;
  (* register *) pwire FA_out_9;
  (* register *) pwire FA_out_10;
  (* register *) pwire FA_out_11;
  (* register *) pwire FA_out_12;
  (* register *) pwire FA_out_13;
  (* register *) pwire FA_out_14;
  (* register *) pwire FA_out_15;
  (* register *) pwire FA_out_16;
  (* register *) pwire FA_out_17;
  (* register *) pwire FA_out_18;
  (* register *) pwire FA_out_19;
  (* register *) pwire FA_out_20;
  (* register *) pwire FA_out_21;
  (* register *) pwire FA_out_22;
  (* register *) pwire FA_out_23;
  (* register *) pwire FA_out_24;
  (* register *) pwire FA_out_25;
  (* register *) pwire FA_out_26;
  (* register *) pwire FA_out_27;
  (* register *) pwire FA_out_28;
  (* register *) pwire FA_out_29;
  (* register *) pwire FA_out_30;
  (* register *) pwire FA_out_31;
  (* register *) pwire FA_out_32;
  (* register *) pwire FA_out_33;
  (* register *) pwire FA_out_34;
  (* register *) pwire FA_out_35;
  (* register *) pwire FA_out_36;
  (* register *) pwire FA_out_37;
  (* register *) pwire FA_out_38;
  (* register *) pwire FA_out_39;
  (* register *) pwire FA_out_40;
  (* register *) pwire FA_out_41;
  (* register *) pwire FA_out_42;
  (* register *) pwire FA_out_43;
  (* register *) pwire FA_out_44;
  (* register *) pwire FA_out_45;
  (* register *) pwire FA_out_46;
  (* register *) pwire FA_out_47;
  (* register *) pwire FA_out_48;
  (* register *) pwire FA_out_49;
  (* register *) pwire FA_out_50;
  (* register *) pwire FA_out_51;
  (* register *) pwire FA_out_52;
  (* register *) pwire FA_out_53;
  (* register *) pwire FA_out_54;
  (* register *) pwire FA_out_55;
  (* register *) pwire FA_out_56;
  (* register *) pwire FA_out_57;
  (* register *) pwire FA_out_58;
  (* register *) pwire FA_out_59;
  (* register *) pwire FA_out_60;
  (* register *) pwire FA_out_61;
  (* register *) pwire FA_out_62;
  (* register *) pwire FA_out_63;
  (* register *) pwire FA_out_64;
  (* register *) pwire FA_out_65;
  (* register *) pwire FA_out_66;
  (* register *) pwire FA_out_67;
  (* register *) pwire FA_out_68;
  (* register *) pwire FA_out_69;
  (* register *) pwire FA_out_70;
  (* register *) pwire FA_out_71;
  (* register *) pwire FA_out_72;
  (* register *) pwire FA_out_73;
  (* register *) pwire FA_out_74;
  (* register *) pwire FA_out_75;
  (* register *) pwire FA_out_76;
  (* register *) pwire FA_out_77;
  (* register *) pwire FA_out_78;
  (* register *) pwire FA_out_79;
  (* register *) pwire FA_out_80;
  (* register *) pwire FA_out_81;
  (* register *) pwire FA_out_82;
  (* register *) pwire FA_out_83;
  (* register *) pwire FA_out_84;
  (* register *) pwire FA_out_85;
  (* register *) pwire FA_out_86;
  (* register *) pwire FA_out_87;
  (* register *) pwire FA_out_88;
  (* register *) pwire FA_out_89;
  (* register *) pwire FA_out_90;
  (* register *) pwire FA_out_91;
  (* register *) pwire FA_out_92;
  (* register *) pwire FA_out_93;
  (* register *) pwire FA_out_94;
  (* register *) pwire FA_out_95;
  (* register *) pwire FA_out_96;
  (* register *) pwire FA_out_97;
  (* register *) pwire FA_out_98;
  (* register *) pwire FA_out_99;
  (* register *) pwire FA_out_100;
  (* register *) pwire FA_out_101;
  (* register *) pwire FA_out_102;
  (* register *) pwire FA_out_103;
  (* register *) pwire FA_out_104;
  (* register *) pwire FA_out_105;
  (* register *) pwire FA_out_106;
  (* register *) pwire FA_out_107;
  (* register *) pwire FA_out_108;
  (* register *) pwire FA_out_109;
  (* register *) pwire FA_out_110;
  (* register *) pwire FA_out_111;
  (* register *) pwire FA_out_112;
  (* register *) pwire FA_out_113;
  (* register *) pwire FA_out_114;
  (* register *) pwire FA_out_115;
  (* register *) pwire FA_out_116;
  (* register *) pwire FA_out_117;
  (* register *) pwire FA_out_118;
  (* register *) pwire FA_out_119;
  (* register *) pwire FA_out_120;
  (* register *) pwire FA_out_121;
  (* register *) pwire FA_out_122;
  (* register *) pwire FA_out_123;
  (* register *) pwire FA_out_124;
  (* register *) pwire FA_out_125;
  (* register *) pwire FA_out_126;
  (* register *) pwire FA_out_127;
  (* register *) pwire FA_out_128;
  (* register *) pwire FA_out_129;
  (* register *) pwire FA_out_130;
  (* register *) pwire FA_out_131;
  (* register *) pwire FA_out_132;
  (* register *) pwire FA_out_133;
  (* register *) pwire FA_out_134;
  (* register *) pwire FA_out_135;
  (* register *) pwire FA_out_136;
  (* register *) pwire FA_out_137;
  (* register *) pwire FA_out_138;
  (* register *) pwire FA_out_139;
  (* register *) pwire FA_out_140;
  (* register *) pwire FA_out_141;
  (* register *) pwire FA_out_142;
  (* register *) pwire FA_out_143;
  (* register *) pwire FA_out_144;
  (* register *) pwire FA_out_145;
  (* register *) pwire FA_out_146;
  (* register *) pwire FA_out_147;
  (* register *) pwire FA_out_148;
  (* register *) pwire FA_out_149;
  (* register *) pwire FA_out_150;
  (* register *) pwire FA_out_151;
  (* register *) pwire FA_out_152;
  (* register *) pwire FA_out_153;
  (* register *) pwire FA_out_154;
  (* register *) pwire FA_out_155;
  (* register *) pwire FA_out_156;
  (* register *) pwire FA_out_157;
  (* register *) pwire FA_out_158;
  (* register *) pwire FA_out_159;
  (* register *) pwire FA_out_160;
  (* register *) pwire FA_out_161;
  (* register *) pwire FA_out_162;
  (* register *) pwire FA_out_163;
  (* register *) pwire FA_out_164;
  (* register *) pwire FA_out_165;
  (* register *) pwire FA_out_166;
  (* register *) pwire FA_out_167;
  (* register *) pwire FA_out_168;
  (* register *) pwire FA_out_169;
  (* register *) pwire FA_out_170;
  (* register *) pwire FA_out_171;
  (* register *) pwire FA_out_172;
  (* register *) pwire FA_out_173;
  (* register *) pwire FA_out_174;
  (* register *) pwire FA_out_175;
  (* register *) pwire FA_out_176;
  (* register *) pwire FA_out_177;
  (* register *) pwire FA_out_178;
  (* register *) pwire FA_out_179;
  (* register *) pwire FA_out_180;
  (* register *) pwire FA_out_181;
  (* register *) pwire FA_out_182;
  (* register *) pwire FA_out_183;
  (* register *) pwire FA_out_184;
  (* register *) pwire FA_out_185;
  (* register *) pwire FA_out_186;
  (* register *) pwire FA_out_187;
  (* register *) pwire FA_out_188;
  (* register *) pwire FA_out_189;
  (* register *) pwire FA_out_190;
  (* register *) pwire FA_out_191;
  (* register *) pwire FA_out_192;
  (* register *) pwire FA_out_193;
  (* register *) pwire FA_out_194;
  (* register *) pwire FA_out_195;
  (* register *) pwire FA_out_196;
  (* register *) pwire FA_out_197;
  (* register *) pwire FA_out_198;
  (* register *) pwire FA_out_199;
  (* register *) pwire FA_out_200;
  (* register *) pwire FA_out_201;
  (* register *) pwire FA_out_202;
  (* register *) pwire FA_out_203;
  (* register *) pwire FA_out_204;
  (* register *) pwire FA_out_205;
  (* register *) pwire FA_out_206;
  (* register *) pwire FA_out_207;
  (* register *) pwire FA_out_208;
  (* register *) pwire FA_out_209;
  (* register *) pwire FA_out_210;
  (* register *) pwire FA_out_211;
  (* register *) pwire FA_out_212;
  (* register *) pwire FA_out_213;
  (* register *) pwire FA_out_214;
  (* register *) pwire FA_out_215;
  (* register *) pwire FA_out_216;
  (* register *) pwire FA_out_217;
  (* register *) pwire FA_out_218;
  (* register *) pwire FA_out_219;
  (* register *) pwire FA_out_220;
  (* register *) pwire FA_out_221;
  (* register *) pwire FA_out_222;
  (* register *) pwire FA_out_223;
  (* register *) pwire FA_out_224;
  (* register *) pwire FA_out_225;
  (* register *) pwire FA_out_226;
  (* register *) pwire FA_out_227;
  (* register *) pwire FA_out_228;
  (* register *) pwire FA_out_229;
  (* register *) pwire FA_out_230;
  (* register *) pwire FA_out_231;
  (* register *) pwire FA_out_232;
  (* register *) pwire FA_out_233;
  (* register *) pwire FA_out_234;
  (* register *) pwire FA_out_235;
  (* register *) pwire FA_out_236;
  (* register *) pwire FA_out_237;
  (* register *) pwire FA_out_238;
  (* register *) pwire FA_out_239;
  (* register *) pwire FA_out_240;
  (* register *) pwire FA_out_241;
  (* register *) pwire FA_out_242;
  (* register *) pwire FA_out_243;
  (* register *) pwire FA_out_244;
  (* register *) pwire FA_out_245;
  (* register *) pwire FA_out_246;
  (* register *) pwire FA_out_247;
  (* register *) pwire FA_out_248;
  (* register *) pwire FA_out_249;
  (* register *) pwire FA_out_250;
  (* register *) pwire FA_out_251;
  (* register *) pwire FA_out_252;
  (* register *) pwire FA_out_253;
  (* register *) pwire FA_out_254;
  (* register *) pwire FA_out_255;
  (* register *) pwire FA_out_256;
  (* register *) pwire FA_out_257;
  (* register *) pwire FA_out_258;
  (* register *) pwire FA_out_259;
  (* register *) pwire FA_out_260;
  (* register *) pwire FA_out_261;
  (* register *) pwire FA_out_262;
  (* register *) pwire FA_out_263;
  (* register *) pwire FA_out_264;
  (* register *) pwire FA_out_265;
  (* register *) pwire FA_out_266;
  (* register *) pwire FA_out_267;
  (* register *) pwire FA_out_268;
  (* register *) pwire FA_out_269;
  (* register *) pwire FA_out_270;
  (* register *) pwire FA_out_271;
  (* register *) pwire FA_out_272;
  (* register *) pwire FA_out_273;
  (* register *) pwire FA_out_274;
  (* register *) pwire FA_out_275;
  (* register *) pwire FA_out_276;
  (* register *) pwire FA_out_277;
  (* register *) pwire FA_out_278;
  (* register *) pwire FA_out_279;
  (* register *) pwire FA_out_280;
  (* register *) pwire FA_out_281;
  (* register *) pwire FA_out_282;
  (* register *) pwire FA_out_283;
  (* register *) pwire FA_out_284;
  (* register *) pwire FA_out_285;
  (* register *) pwire FA_out_286;
  (* register *) pwire FA_out_287;
  (* register *) pwire FA_out_288;
  (* register *) pwire FA_out_289;
  (* register *) pwire FA_out_290;
  (* register *) pwire FA_out_291;
  (* register *) pwire FA_out_292;
  (* register *) pwire FA_out_293;
  (* register *) pwire FA_out_294;
  (* register *) pwire FA_out_295;
  (* register *) pwire FA_out_296;
  (* register *) pwire FA_out_297;
  (* register *) pwire FA_out_298;
  (* register *) pwire FA_out_299;
  (* register *) pwire FA_out_300;
  (* register *) pwire FA_out_301;
  (* register *) pwire FA_out_302;
  (* register *) pwire FA_out_303;
  (* register *) pwire FA_out_304;
  (* register *) pwire FA_out_305;
  (* register *) pwire FA_out_306;
  (* register *) pwire FA_out_307;
  (* register *) pwire FA_out_308;
  (* register *) pwire FA_out_309;
  (* register *) pwire FA_out_310;
  (* register *) pwire FA_out_311;
  (* register *) pwire FA_out_312;
  (* register *) pwire FA_out_313;
  (* register *) pwire FA_out_314;
  (* register *) pwire FA_out_315;
  (* register *) pwire FA_out_316;
  (* register *) pwire FA_out_317;
  (* register *) pwire FA_out_318;
  (* register *) pwire FA_out_319;
  (* register *) pwire FA_out_320;
  (* register *) pwire FA_out_321;
  (* register *) pwire FA_out_322;
  (* register *) pwire FA_out_323;
  (* register *) pwire FA_out_324;
  (* register *) pwire FA_out_325;
  (* register *) pwire FA_out_326;
  (* register *) pwire FA_out_327;
  (* register *) pwire FA_out_328;
  (* register *) pwire FA_out_329;
  (* register *) pwire FA_out_330;
  (* register *) pwire FA_out_331;
  (* register *) pwire FA_out_332;
  (* register *) pwire FA_out_333;
  (* register *) pwire FA_out_334;
  (* register *) pwire FA_out_335;
  (* register *) pwire FA_out_336;
  (* register *) pwire FA_out_337;
  (* register *) pwire FA_out_338;
  (* register *) pwire FA_out_339;
  (* register *) pwire FA_out_340;
  (* register *) pwire FA_out_341;
  (* register *) pwire FA_out_342;
  (* register *) pwire FA_out_343;
  (* register *) pwire FA_out_344;
  (* register *) pwire FA_out_345;
  (* register *) pwire FA_out_346;
  (* register *) pwire FA_out_347;
  (* register *) pwire FA_out_348;
  (* register *) pwire FA_out_349;
  (* register *) pwire FA_out_350;
  (* register *) pwire FA_out_351;
  (* register *) pwire FA_out_352;
  (* register *) pwire FA_out_353;
  (* register *) pwire FA_out_354;
  (* register *) pwire FA_out_355;
  (* register *) pwire FA_out_356;
  (* register *) pwire FA_out_357;
  (* register *) pwire FA_out_358;
  (* register *) pwire FA_out_359;
  (* register *) pwire FA_out_360;
  (* register *) pwire FA_out_361;
  (* register *) pwire FA_out_362;
  (* register *) pwire FA_out_363;
  (* register *) pwire FA_out_364;
  (* register *) pwire FA_out_365;
  (* register *) pwire FA_out_366;
  (* register *) pwire FA_out_367;
  (* register *) pwire FA_out_368;
  (* register *) pwire FA_out_369;
  (* register *) pwire FA_out_370;
  (* register *) pwire FA_out_371;
  (* register *) pwire FA_out_372;
  (* register *) pwire FA_out_373;
  (* register *) pwire FA_out_374;
  (* register *) pwire FA_out_375;
  (* register *) pwire FA_out_376;
  (* register *) pwire FA_out_377;
  (* register *) pwire FA_out_378;
  (* register *) pwire FA_out_379;
  (* register *) pwire FA_out_380;
  (* register *) pwire FA_out_381;
  (* register *) pwire FA_out_382;
  (* register *) pwire FA_out_383;
  (* register *) pwire FA_out_384;
  (* register *) pwire FA_out_385;
  (* register *) pwire FA_out_386;
  (* register *) pwire FA_out_387;
  (* register *) pwire FA_out_388;
  (* register *) pwire FA_out_389;
  (* register *) pwire FA_out_390;
  (* register *) pwire FA_out_391;
  (* register *) pwire FA_out_392;
  (* register *) pwire FA_out_393;
  (* register *) pwire FA_out_394;
  (* register *) pwire FA_out_395;
  (* register *) pwire FA_out_396;
  (* register *) pwire FA_out_397;
  (* register *) pwire FA_out_398;
  (* register *) pwire FA_out_399;
  (* register *) pwire FA_out_400;
  (* register *) pwire FA_out_401;
  (* register *) pwire FA_out_402;
  (* register *) pwire FA_out_403;
  (* register *) pwire FA_out_404;
  (* register *) pwire FA_out_405;
  (* register *) pwire FA_out_406;
  (* register *) pwire FA_out_407;
  (* register *) pwire FA_out_408;
  (* register *) pwire FA_out_409;
  (* register *) pwire FA_out_410;
  (* register *) pwire FA_out_411;
  (* register *) pwire FA_out_412;
  (* register *) pwire FA_out_413;
  (* register *) pwire FA_out_414;
  (* register *) pwire FA_out_415;
  (* register *) pwire FA_out_416;
  (* register *) pwire FA_out_417;
  (* register *) pwire FA_out_418;
  (* register *) pwire FA_out_419;
  (* register *) pwire FA_out_420;
  (* register *) pwire FA_out_421;
  (* register *) pwire FA_out_422;
  (* register *) pwire FA_out_423;
  (* register *) pwire FA_out_424;
  (* register *) pwire FA_out_425;
  (* register *) pwire FA_out_426;
  (* register *) pwire FA_out_427;
  (* register *) pwire FA_out_428;
  (* register *) pwire FA_out_429;
  (* register *) pwire FA_out_430;
  (* register *) pwire FA_out_431;
  (* register *) pwire FA_out_432;
  (* register *) pwire FA_out_433;
  (* register *) pwire FA_out_434;
  (* register *) pwire FA_out_435;
  (* register *) pwire FA_out_436;
  (* register *) pwire FA_out_437;
  (* register *) pwire FA_out_438;
  (* register *) pwire FA_out_439;
  (* register *) pwire FA_out_440;
  (* register *) pwire FA_out_441;
  (* register *) pwire FA_out_442;
  (* register *) pwire FA_out_443;
  (* register *) pwire FA_out_444;
  (* register *) pwire FA_out_445;
  (* register *) pwire FA_out_446;
  (* register *) pwire FA_out_447;
  (* register *) pwire FA_out_448;
  (* register *) pwire FA_out_449;
  (* register *) pwire FA_out_450;
  (* register *) pwire FA_out_451;
  (* register *) pwire FA_out_452;
  (* register *) pwire FA_out_453;
  (* register *) pwire FA_out_454;
  (* register *) pwire FA_out_455;
  (* register *) pwire FA_out_456;
  (* register *) pwire FA_out_457;
  (* register *) pwire FA_out_458;
  (* register *) pwire FA_out_459;
  (* register *) pwire FA_out_460;
  (* register *) pwire FA_out_461;
  (* register *) pwire FA_out_462;
  (* register *) pwire FA_out_463;
  (* register *) pwire FA_out_464;
  (* register *) pwire FA_out_465;
  (* register *) pwire FA_out_466;
  (* register *) pwire FA_out_467;
  (* register *) pwire FA_out_468;
  (* register *) pwire FA_out_469;
  (* register *) pwire FA_out_470;
  (* register *) pwire FA_out_471;
  (* register *) pwire FA_out_472;
  (* register *) pwire FA_out_473;
  (* register *) pwire FA_out_474;
  (* register *) pwire FA_out_475;
  (* register *) pwire FA_out_476;
  (* register *) pwire FA_out_477;
  (* register *) pwire FA_out_478;
  (* register *) pwire FA_out_479;
  (* register *) pwire FA_out_480;
  (* register *) pwire FA_out_481;
  (* register *) pwire FA_out_482;
  (* register *) pwire FA_out_483;
  (* register *) pwire FA_out_484;
  (* register *) pwire FA_out_485;
  (* register *) pwire FA_out_486;
  (* register *) pwire FA_out_487;
  (* register *) pwire FA_out_488;
  (* register *) pwire FA_out_489;
  (* register *) pwire FA_out_490;
  (* register *) pwire FA_out_491;
  (* register *) pwire FA_out_492;
  (* register *) pwire FA_out_493;
  (* register *) pwire FA_out_494;
  (* register *) pwire FA_out_495;
  (* register *) pwire FA_out_496;
  (* register *) pwire FA_out_497;
  (* register *) pwire FA_out_498;
  (* register *) pwire FA_out_499;
  (* register *) pwire FA_out_500;
  (* register *) pwire FA_out_501;
  (* register *) pwire FA_out_502;
  (* register *) pwire FA_out_503;
  (* register *) pwire FA_out_504;
  (* register *) pwire FA_out_505;
  (* register *) pwire FA_out_506;
  (* register *) pwire FA_out_507;
  (* register *) pwire FA_out_508;
  (* register *) pwire FA_out_509;
  (* register *) pwire FA_out_510;
  (* register *) pwire FA_out_511;
  (* register *) pwire FA_out_512;
  (* register *) pwire FA_out_513;
  (* register *) pwire FA_out_514;
  (* register *) pwire FA_out_515;
  (* register *) pwire FA_out_516;
  (* register *) pwire FA_out_517;
  (* register *) pwire FA_out_518;
  (* register *) pwire FA_out_519;
  (* register *) pwire FA_out_520;
  (* register *) pwire FA_out_521;
  (* register *) pwire FA_out_522;
  (* register *) pwire FA_out_523;
  (* register *) pwire FA_out_524;
  (* register *) pwire FA_out_525;
  (* register *) pwire FA_out_526;
  (* register *) pwire FA_out_527;
  (* register *) pwire FA_out_528;
  (* register *) pwire FA_out_529;
  (* register *) pwire FA_out_530;
  (* register *) pwire FA_out_531;
  (* register *) pwire FA_out_532;
  (* register *) pwire FA_out_533;
  (* register *) pwire FA_out_534;
  (* register *) pwire FA_out_535;
  (* register *) pwire FA_out_536;
  (* register *) pwire FA_out_537;
  (* register *) pwire FA_out_538;
  (* register *) pwire FA_out_539;
  (* register *) pwire FA_out_540;
  (* register *) pwire FA_out_541;
  (* register *) pwire FA_out_542;
  (* register *) pwire FA_out_543;
  (* register *) pwire FA_out_544;
  (* register *) pwire FA_out_545;
  (* register *) pwire FA_out_546;
  (* register *) pwire FA_out_547;
  (* register *) pwire FA_out_548;
  (* register *) pwire FA_out_549;
  (* register *) pwire FA_out_550;
  (* register *) pwire FA_out_551;
  (* register *) pwire FA_out_552;
  (* register *) pwire FA_out_553;
  (* register *) pwire FA_out_554;
  (* register *) pwire FA_out_555;
  (* register *) pwire FA_out_556;
  (* register *) pwire FA_out_557;
  (* register *) pwire FA_out_558;
  (* register *) pwire FA_out_559;
  (* register *) pwire FA_out_560;
  (* register *) pwire FA_out_561;
  (* register *) pwire FA_out_562;
  (* register *) pwire FA_out_563;
  (* register *) pwire FA_out_564;
  (* register *) pwire FA_out_565;
  (* register *) pwire FA_out_566;
  (* register *) pwire FA_out_567;
  (* register *) pwire FA_out_568;
  (* register *) pwire FA_out_569;
  (* register *) pwire FA_out_570;
  (* register *) pwire FA_out_571;
  (* register *) pwire FA_out_572;
  (* register *) pwire FA_out_573;
  (* register *) pwire FA_out_574;
  (* register *) pwire FA_out_575;
  (* register *) pwire FA_out_576;
  (* register *) pwire FA_out_577;
  (* register *) pwire FA_out_578;
  (* register *) pwire FA_out_579;
  (* register *) pwire FA_out_580;
  (* register *) pwire FA_out_581;
  (* register *) pwire FA_out_582;
  (* register *) pwire FA_out_583;
  (* register *) pwire FA_out_584;
  (* register *) pwire FA_out_585;
  (* register *) pwire FA_out_586;
  (* register *) pwire FA_out_587;
  (* register *) pwire FA_out_588;
  (* register *) pwire FA_out_589;
  (* register *) pwire FA_out_590;
  (* register *) pwire FA_out_591;
  (* register *) pwire FA_out_592;
  (* register *) pwire FA_out_593;
  (* register *) pwire FA_out_594;
  (* register *) pwire FA_out_595;
  (* register *) pwire FA_out_596;
  (* register *) pwire FA_out_597;
  (* register *) pwire FA_out_598;
  (* register *) pwire FA_out_599;
  (* register *) pwire FA_out_600;
  (* register *) pwire FA_out_601;
  (* register *) pwire FA_out_602;
  (* register *) pwire FA_out_603;
  (* register *) pwire FA_out_604;
  (* register *) pwire FA_out_605;
  (* register *) pwire FA_out_606;
  (* register *) pwire FA_out_607;
  (* register *) pwire FA_out_608;
  (* register *) pwire FA_out_609;
  (* register *) pwire FA_out_610;
  (* register *) pwire FA_out_611;
  (* register *) pwire FA_out_612;
  (* register *) pwire FA_out_613;
  (* register *) pwire FA_out_614;
  (* register *) pwire FA_out_615;
  (* register *) pwire FA_out_616;
  (* register *) pwire FA_out_617;
  (* register *) pwire FA_out_618;
  (* register *) pwire FA_out_619;
  (* register *) pwire FA_out_620;
  (* register *) pwire FA_out_621;
  (* register *) pwire FA_out_622;
  (* register *) pwire FA_out_623;
  (* register *) pwire FA_out_624;
  (* register *) pwire FA_out_625;
  (* register *) pwire FA_out_626;
  (* register *) pwire FA_out_627;
  (* register *) pwire FA_out_628;
  (* register *) pwire FA_out_629;
  (* register *) pwire FA_out_630;
  (* register *) pwire FA_out_631;
  (* register *) pwire FA_out_632;
  (* register *) pwire FA_out_633;
  (* register *) pwire FA_out_634;
  (* register *) pwire FA_out_635;
  (* register *) pwire FA_out_636;
  (* register *) pwire FA_out_637;
  (* register *) pwire FA_out_638;
  (* register *) pwire FA_out_639;
  (* register *) pwire FA_out_640;
  (* register *) pwire FA_out_641;
  (* register *) pwire FA_out_642;
  (* register *) pwire FA_out_643;
  (* register *) pwire FA_out_644;
  (* register *) pwire FA_out_645;
  (* register *) pwire FA_out_646;
  (* register *) pwire FA_out_647;
  (* register *) pwire FA_out_648;
  (* register *) pwire FA_out_649;
  (* register *) pwire FA_out_650;
  (* register *) pwire FA_out_651;
  (* register *) pwire FA_out_652;
  (* register *) pwire FA_out_653;
  (* register *) pwire FA_out_654;
  (* register *) pwire FA_out_655;
  (* register *) pwire FA_out_656;
  (* register *) pwire FA_out_657;
  (* register *) pwire FA_out_658;
  (* register *) pwire FA_out_659;
  (* register *) pwire FA_out_660;
  (* register *) pwire FA_out_661;
  (* register *) pwire FA_out_662;
  (* register *) pwire FA_out_663;
  (* register *) pwire FA_out_664;
  (* register *) pwire FA_out_665;
  (* register *) pwire FA_out_666;
  (* register *) pwire FA_out_667;
  (* register *) pwire FA_out_668;
  (* register *) pwire FA_out_669;
  (* register *) pwire FA_out_670;
  (* register *) pwire FA_out_671;
  (* register *) pwire FA_out_672;
  (* register *) pwire FA_out_673;
  (* register *) pwire FA_out_674;
  (* register *) pwire FA_out_675;
  (* register *) pwire FA_out_676;
  (* register *) pwire FA_out_677;
  (* register *) pwire FA_out_678;
  (* register *) pwire FA_out_679;
  (* register *) pwire FA_out_680;
  (* register *) pwire FA_out_681;
  (* register *) pwire FA_out_682;
  (* register *) pwire FA_out_683;
  (* register *) pwire FA_out_684;
  (* register *) pwire FA_out_685;
  (* register *) pwire FA_out_686;
  (* register *) pwire FA_out_687;
  (* register *) pwire FA_out_688;
  (* register *) pwire FA_out_689;
  (* register *) pwire FA_out_690;
  (* register *) pwire FA_out_691;
  (* register *) pwire FA_out_692;
  (* register *) pwire FA_out_693;
  (* register *) pwire FA_out_694;
  (* register *) pwire FA_out_695;
  (* register *) pwire FA_out_696;
  (* register *) pwire FA_out_697;
  (* register *) pwire FA_out_698;
  (* register *) pwire FA_out_699;
  (* register *) pwire FA_out_700;
  (* register *) pwire FA_out_701;
  (* register *) pwire FA_out_702;
  (* register *) pwire FA_out_703;
  (* register *) pwire FA_out_704;
  (* register *) pwire FA_out_705;
  (* register *) pwire FA_out_706;
  (* register *) pwire FA_out_707;
  (* register *) pwire FA_out_708;
  (* register *) pwire FA_out_709;
  (* register *) pwire FA_out_710;
  (* register *) pwire FA_out_711;
  (* register *) pwire FA_out_712;
  (* register *) pwire FA_out_713;
  (* register *) pwire FA_out_714;
  (* register *) pwire FA_out_715;
  (* register *) pwire FA_out_716;
  (* register *) pwire FA_out_717;
  (* register *) pwire FA_out_718;
  (* register *) pwire FA_out_719;
  (* register *) pwire FA_out_720;
  (* register *) pwire FA_out_721;
  (* register *) pwire FA_out_722;
  (* register *) pwire FA_out_723;
  (* register *) pwire FA_out_724;
  (* register *) pwire FA_out_725;
  (* register *) pwire FA_out_726;
  (* register *) pwire FA_out_727;
  (* register *) pwire FA_out_728;
  (* register *) pwire FA_out_729;
  (* register *) pwire FA_out_730;
  (* register *) pwire FA_out_731;
  (* register *) pwire FA_out_732;
  (* register *) pwire FA_out_733;
  (* register *) pwire FA_out_734;
  (* register *) pwire FA_out_735;
  (* register *) pwire FA_out_736;
  (* register *) pwire FA_out_737;
  (* register *) pwire FA_out_738;
  (* register *) pwire FA_out_739;
  (* register *) pwire FA_out_740;
  (* register *) pwire FA_out_741;
  (* register *) pwire FA_out_742;
  (* register *) pwire FA_out_743;
  (* register *) pwire FA_out_744;
  (* register *) pwire FA_out_745;
  (* register *) pwire FA_out_746;
  (* register *) pwire FA_out_747;
  (* register *) pwire FA_out_748;
  (* register *) pwire FA_out_749;
  (* register *) pwire FA_out_750;
  (* register *) pwire FA_out_751;
  (* register *) pwire FA_out_752;
  (* register *) pwire FA_out_753;
  (* register *) pwire FA_out_754;
  (* register *) pwire FA_out_755;
  (* register *) pwire FA_out_756;
  (* register *) pwire FA_out_757;
  (* register *) pwire FA_out_758;
  (* register *) pwire FA_out_759;
  (* register *) pwire FA_out_760;
  (* register *) pwire FA_out_761;
  (* register *) pwire FA_out_762;
  (* register *) pwire FA_out_763;
  (* register *) pwire FA_out_764;
  (* register *) pwire FA_out_765;
  (* register *) pwire FA_out_766;
  (* register *) pwire FA_out_767;
  (* register *) pwire FA_out_768;
  (* register *) pwire FA_out_769;
  (* register *) pwire FA_out_770;
  (* register *) pwire FA_out_771;
  (* register *) pwire FA_out_772;
  (* register *) pwire FA_out_773;
  (* register *) pwire FA_out_774;
  (* register *) pwire FA_out_775;
  (* register *) pwire FA_out_776;
  (* register *) pwire FA_out_777;
  (* register *) pwire FA_out_778;
  (* register *) pwire FA_out_779;
  (* register *) pwire FA_out_780;
  (* register *) pwire FA_out_781;
  (* register *) pwire FA_out_782;
  (* register *) pwire FA_out_783;
  (* register *) pwire FA_out_784;
  (* register *) pwire FA_out_785;
  (* register *) pwire FA_out_786;
  (* register *) pwire FA_out_787;
  (* register *) pwire FA_out_788;
  (* register *) pwire FA_out_789;
  (* register *) pwire FA_out_790;
  (* register *) pwire FA_out_791;
  (* register *) pwire FA_out_792;
  (* register *) pwire FA_out_793;
  (* register *) pwire FA_out_794;
  (* register *) pwire FA_out_795;
  (* register *) pwire FA_out_796;
  (* register *) pwire FA_out_797;
  (* register *) pwire FA_out_798;
  (* register *) pwire FA_out_799;
  (* register *) pwire FA_out_800;
  (* register *) pwire FA_out_801;
  (* register *) pwire FA_out_802;
  (* register *) pwire FA_out_803;
  (* register *) pwire FA_out_804;
  (* register *) pwire FA_out_805;
  (* register *) pwire FA_out_806;
  (* register *) pwire FA_out_807;
  (* register *) pwire FA_out_808;
  (* register *) pwire FA_out_809;
  (* register *) pwire FA_out_810;
  (* register *) pwire FA_out_811;
  (* register *) pwire FA_out_812;
  (* register *) pwire FA_out_813;
  (* register *) pwire FA_out_814;
  (* register *) pwire FA_out_815;
  (* register *) pwire FA_out_816;
  (* register *) pwire FA_out_817;
  (* register *) pwire FA_out_818;
  (* register *) pwire FA_out_819;
  (* register *) pwire FA_out_820;
  (* register *) pwire FA_out_821;
  (* register *) pwire FA_out_822;
  (* register *) pwire FA_out_823;
  (* register *) pwire FA_out_824;
  (* register *) pwire FA_out_825;
  (* register *) pwire FA_out_826;
  (* register *) pwire FA_out_827;
  (* register *) pwire FA_out_828;
  (* register *) pwire FA_out_829;
  (* register *) pwire FA_out_830;
  (* register *) pwire FA_out_831;
  (* register *) pwire FA_out_832;
  (* register *) pwire FA_out_833;
  (* register *) pwire FA_out_834;
  (* register *) pwire FA_out_835;
  (* register *) pwire FA_out_836;
  (* register *) pwire FA_out_837;
  (* register *) pwire FA_out_838;
  (* register *) pwire FA_out_839;
  (* register *) pwire FA_out_840;
  (* register *) pwire FA_out_841;
  (* register *) pwire FA_out_842;
  (* register *) pwire FA_out_843;
  (* register *) pwire FA_out_844;
  (* register *) pwire FA_out_845;
  (* register *) pwire FA_out_846;
  (* register *) pwire FA_out_847;
  (* register *) pwire FA_out_848;
  (* register *) pwire FA_out_849;
  (* register *) pwire FA_out_850;
  (* register *) pwire FA_out_851;
  (* register *) pwire FA_out_852;
  (* register *) pwire FA_out_853;
  (* register *) pwire FA_out_854;
  (* register *) pwire FA_out_855;
  (* register *) pwire FA_out_856;
  (* register *) pwire FA_out_857;
  (* register *) pwire FA_out_858;
  (* register *) pwire FA_out_859;
  (* register *) pwire FA_out_860;
  (* register *) pwire FA_out_861;
  (* register *) pwire FA_out_862;
  (* register *) pwire FA_out_863;
  (* register *) pwire FA_out_864;
  (* register *) pwire FA_out_865;
  (* register *) pwire FA_out_866;
  (* register *) pwire FA_out_867;
  (* register *) pwire FA_out_868;
  (* register *) pwire FA_out_869;
  (* register *) pwire FA_out_870;
  (* register *) pwire FA_out_871;
  (* register *) pwire FA_out_872;
  (* register *) pwire FA_out_873;
  (* register *) pwire FA_out_874;
  (* register *) pwire FA_out_875;
  (* register *) pwire FA_out_876;
  (* register *) pwire FA_out_877;
  (* register *) pwire FA_out_878;
  (* register *) pwire FA_out_879;
  (* register *) pwire FA_out_880;
  (* register *) pwire FA_out_881;
  (* register *) pwire FA_out_882;
  (* register *) pwire FA_out_883;
  (* register *) pwire FA_out_884;
  (* register *) pwire FA_out_885;
  (* register *) pwire FA_out_886;
  (* register *) pwire FA_out_887;
  (* register *) pwire FA_out_888;
  (* register *) pwire FA_out_889;
  (* register *) pwire FA_out_890;
  (* register *) pwire FA_out_891;
  (* register *) pwire FA_out_892;
  (* register *) pwire FA_out_893;
  (* register *) pwire FA_out_894;
  (* register *) pwire FA_out_895;
  (* register *) pwire FA_out_896;
  (* register *) pwire FA_out_897;
  (* register *) pwire FA_out_898;
  (* register *) pwire FA_out_899;
  (* register *) pwire FA_out_900;
  (* register *) pwire FA_out_901;
  (* register *) pwire FA_out_902;
  (* register *) pwire FA_out_903;
  (* register *) pwire FA_out_904;
  (* register *) pwire FA_out_905;
  (* register *) pwire FA_out_906;
  (* register *) pwire FA_out_907;
  (* register *) pwire FA_out_908;
  (* register *) pwire FA_out_909;
  (* register *) pwire FA_out_910;
  (* register *) pwire FA_out_911;
  (* register *) pwire FA_out_912;
  (* register *) pwire FA_out_913;
  (* register *) pwire FA_out_914;
  (* register *) pwire FA_out_915;
  (* register *) pwire FA_out_916;
  (* register *) pwire FA_out_917;
  (* register *) pwire FA_out_918;
  (* register *) pwire FA_out_919;
  (* register *) pwire FA_out_920;
  (* register *) pwire FA_out_921;
  (* register *) pwire FA_out_922;
  (* register *) pwire FA_out_923;
  (* register *) pwire FA_out_924;
  (* register *) pwire FA_out_925;
  (* register *) pwire FA_out_926;
  (* register *) pwire FA_out_927;
  (* register *) pwire FA_out_928;
  (* register *) pwire FA_out_929;
  (* register *) pwire FA_out_930;
  (* register *) pwire FA_out_931;
  (* register *) pwire FA_out_932;
  (* register *) pwire FA_out_933;
  (* register *) pwire FA_out_934;
  (* register *) pwire FA_out_935;
  (* register *) pwire FA_out_936;
  (* register *) pwire FA_out_937;
  (* register *) pwire FA_out_938;
  (* register *) pwire FA_out_939;
  (* register *) pwire FA_out_940;
  (* register *) pwire FA_out_941;
  (* register *) pwire FA_out_942;
  (* register *) pwire FA_out_943;
  (* register *) pwire FA_out_944;
  (* register *) pwire FA_out_945;
  (* register *) pwire FA_out_946;
  (* register *) pwire FA_out_947;
  (* register *) pwire FA_out_948;
  (* register *) pwire FA_out_949;
  (* register *) pwire FA_out_950;
  (* register *) pwire FA_out_951;
  (* register *) pwire FA_out_952;
  (* register *) pwire FA_out_953;
  (* register *) pwire FA_out_954;
  (* register *) pwire FA_out_955;
  (* register *) pwire FA_out_956;
  (* register *) pwire FA_out_957;
  (* register *) pwire FA_out_958;
  (* register *) pwire FA_out_959;
  (* register *) pwire FA_out_960;
  (* register *) pwire FA_out_961;
  (* register *) pwire FA_out_962;
  (* register *) pwire FA_out_963;
  (* register *) pwire FA_out_964;
  (* register *) pwire FA_out_965;
  (* register *) pwire FA_out_966;
  (* register *) pwire FA_out_967;
  (* register *) pwire FA_out_968;
  (* register *) pwire FA_out_969;
  (* register *) pwire FA_out_970;
  (* register *) pwire FA_out_971;
  (* register *) pwire FA_out_972;
  (* register *) pwire FA_out_973;
  (* register *) pwire FA_out_974;
  (* register *) pwire FA_out_975;
  (* register *) pwire FA_out_976;
  (* register *) pwire FA_out_977;
  (* register *) pwire FA_out_978;
  (* register *) pwire FA_out_979;
  (* register *) pwire FA_out_980;
  (* register *) pwire FA_out_981;
  (* register *) pwire FA_out_982;
  (* register *) pwire FA_out_983;
  (* register *) pwire FA_out_984;
  (* register *) pwire FA_out_985;
  (* register *) pwire FA_out_986;
  (* register *) pwire FA_out_987;
  (* register *) pwire FA_out_988;
  (* register *) pwire FA_out_989;
  (* register *) pwire FA_out_990;
  (* register *) pwire FA_out_991;
  (* register *) pwire FA_out_992;
  (* register *) pwire FA_out_993;
  (* register *) pwire FA_out_994;
  (* register *) pwire FA_out_995;
  (* register *) pwire FA_out_996;
  (* register *) pwire FA_out_997;
  (* register *) pwire FA_out_998;
  (* register *) pwire FA_out_999;
  (* register *) pwire FA_out_1000;
  (* register *) pwire FA_out_1001;
  (* register *) pwire FA_out_1002;
  (* register *) pwire FA_out_1003;
  (* register *) pwire FA_out_1004;
  (* register *) pwire FA_out_1005;
  (* register *) pwire FA_out_1006;
  (* register *) pwire FA_out_1007;
  (* register *) pwire FA_out_1008;
  (* register *) pwire FA_out_1009;
  (* register *) pwire FA_out_1010;
  (* register *) pwire FA_out_1011;
  (* register *) pwire FA_out_1012;
  (* register *) pwire FA_out_1013;
  (* register *) pwire FA_out_1014;
  (* register *) pwire FA_out_1015;
  (* register *) pwire FA_out_1016;
  (* register *) pwire FA_out_1017;
  (* register *) pwire FA_out_1018;
  (* register *) pwire FA_out_1019;
  (* register *) pwire FA_out_1020;
  (* register *) pwire FA_out_1021;
  (* register *) pwire FA_out_1022;
  (* register *) pwire FA_out_1023;
  (* register *) pwire FA_out_1024;
  (* register *) pwire FA_out_1025;
  (* register *) pwire FA_out_1026;
  (* register *) pwire FA_out_1027;
  (* register *) pwire FA_out_1028;
  (* register *) pwire FA_out_1029;
  (* register *) pwire FA_out_1030;
  (* register *) pwire FA_out_1031;
  (* register *) pwire FA_out_1032;
  (* register *) pwire FA_out_1033;
  (* register *) pwire FA_out_1034;
  (* register *) pwire FA_out_1035;
  (* register *) pwire FA_out_1036;
  (* register *) pwire FA_out_1037;
  (* register *) pwire FA_out_1038;
  (* register *) pwire FA_out_1039;
  (* register *) pwire FA_out_1040;
  (* register *) pwire FA_out_1041;
  (* register *) pwire FA_out_1042;
  (* register *) pwire FA_out_1043;
  (* register *) pwire FA_out_1044;
  (* register *) pwire FA_out_1045;
  (* register *) pwire FA_out_1046;
  (* register *) pwire FA_out_1047;
  (* register *) pwire FA_out_1048;
  (* register *) pwire FA_out_1049;
  (* register *) pwire FA_out_1050;
  (* register *) pwire FA_out_1051;
  (* register *) pwire FA_out_1052;
  (* register *) pwire FA_out_1053;
  (* register *) pwire FA_out_1054;
  (* register *) pwire FA_out_1055;
  (* register *) pwire FA_out_1056;
  (* register *) pwire FA_out_1057;
  (* register *) pwire FA_out_1058;
  (* register *) pwire FA_out_1059;
  (* register *) pwire FA_out_1060;
  (* register *) pwire FA_out_1061;
  (* register *) pwire FA_out_1062;
  (* register *) pwire FA_out_1063;
  (* register *) pwire FA_out_1064;
  (* register *) pwire FA_out_1065;
  (* register *) pwire FA_out_1066;
  (* register *) pwire FA_out_1067;
  (* register *) pwire FA_out_1068;
  (* register *) pwire FA_out_1069;
  (* register *) pwire FA_out_1070;
  (* register *) pwire FA_out_1071;
  (* register *) pwire FA_out_1072;
  (* register *) pwire FA_out_1073;
  (* register *) pwire FA_out_1074;
  (* register *) pwire FA_out_1075;
  (* register *) pwire FA_out_1076;
  (* register *) pwire FA_out_1077;
  (* register *) pwire FA_out_1078;
  (* register *) pwire FA_out_1079;
  (* register *) pwire FA_out_1080;
  (* register *) pwire FA_out_1081;
  (* register *) pwire FA_out_1082;
  (* register *) pwire FA_out_1083;
  (* register *) pwire FA_out_1084;
  (* register *) pwire FA_out_1085;
  (* register *) pwire FA_out_1086;
  (* register *) pwire FA_out_1087;
  (* register *) pwire FA_out_1088;
  (* register *) pwire FA_out_1089;
  (* register *) pwire FA_out_1090;
  (* register *) pwire FA_out_1091;
  (* register *) pwire FA_out_1092;
  (* register *) pwire FA_out_1093;
  (* register *) pwire FA_out_1094;
  (* register *) pwire FA_out_1095;
  (* register *) pwire FA_out_1096;
  (* register *) pwire FA_out_1097;
  (* register *) pwire FA_out_1098;
  (* register *) pwire FA_out_1099;
  (* register *) pwire FA_out_1100;
  (* register *) pwire FA_out_1101;
  (* register *) pwire FA_out_1102;
  (* register *) pwire FA_out_1103;
  (* register *) pwire FA_out_1104;
  (* register *) pwire FA_out_1105;
  (* register *) pwire FA_out_1106;
  (* register *) pwire FA_out_1107;
  (* register *) pwire FA_out_1108;
  (* register *) pwire FA_out_1109;
  (* register *) pwire FA_out_1110;
  (* register *) pwire FA_out_1111;
  (* register *) pwire FA_out_1112;
  (* register *) pwire FA_out_1113;
  (* register *) pwire FA_out_1114;
  (* register *) pwire FA_out_1115;
  (* register *) pwire FA_out_1116;
  (* register *) pwire FA_out_1117;
  (* register *) pwire FA_out_1118;
  (* register *) pwire FA_out_1119;
  (* register *) pwire FA_out_1120;
  (* register *) pwire FA_out_1121;
  (* register *) pwire FA_out_1122;
  (* register *) pwire FA_out_1123;
  (* register *) pwire FA_out_1124;
  (* register *) pwire FA_out_1125;
  (* register *) pwire FA_out_1126;
  (* register *) pwire FA_out_1127;
  (* register *) pwire FA_out_1128;
  (* register *) pwire FA_out_1129;
  (* register *) pwire FA_out_1130;
  (* register *) pwire FA_out_1131;
  (* register *) pwire FA_out_1132;
  (* register *) pwire FA_out_1133;
  (* register *) pwire FA_out_1134;
  (* register *) pwire FA_out_1135;
  (* register *) pwire FA_out_1136;
  (* register *) pwire FA_out_1137;
  (* register *) pwire FA_out_1138;
  (* register *) pwire FA_out_1139;
  (* register *) pwire FA_out_1140;
  (* register *) pwire FA_out_1141;
  (* register *) pwire FA_out_1142;
  (* register *) pwire FA_out_1143;
  (* register *) pwire FA_out_1144;
  (* register *) pwire FA_out_1145;
  (* register *) pwire FA_out_1146;
  (* register *) pwire FA_out_1147;
  (* register *) pwire FA_out_1148;
  (* register *) pwire FA_out_1149;
  (* register *) pwire FA_out_1150;
  (* register *) pwire FA_out_1151;
  (* register *) pwire FA_out_1152;
  (* register *) pwire FA_out_1153;
  (* register *) pwire FA_out_1154;
  (* register *) pwire FA_out_1155;
  (* register *) pwire FA_out_1156;
  (* register *) pwire FA_out_1157;
  (* register *) pwire FA_out_1158;
  (* register *) pwire FA_out_1159;
  (* register *) pwire FA_out_1160;
  (* register *) pwire FA_out_1161;
  (* register *) pwire FA_out_1162;
  (* register *) pwire FA_out_1163;
  (* register *) pwire FA_out_1164;
  (* register *) pwire FA_out_1165;
  (* register *) pwire FA_out_1166;
  (* register *) pwire FA_out_1167;
  (* register *) pwire FA_out_1168;
  (* register *) pwire FA_out_1169;
  (* register *) pwire FA_out_1170;
  (* register *) pwire FA_out_1171;
  (* register *) pwire FA_out_1172;
  (* register *) pwire FA_out_1173;
  (* register *) pwire FA_out_1174;
  (* register *) pwire FA_out_1175;
  (* register *) pwire FA_out_1176;
  (* register *) pwire FA_out_1177;
  (* register *) pwire FA_out_1178;
  (* register *) pwire FA_out_1179;
  (* register *) pwire FA_out_1180;
  (* register *) pwire FA_out_1181;
  (* register *) pwire FA_out_1182;
  (* register *) pwire FA_out_1183;
  (* register *) pwire FA_out_1184;
  (* register *) pwire FA_out_1185;
  (* register *) pwire FA_out_1186;
  (* register *) pwire FA_out_1187;
  (* register *) pwire FA_out_1188;
  (* register *) pwire FA_out_1189;
  (* register *) pwire FA_out_1190;
  (* register *) pwire FA_out_1191;
  (* register *) pwire FA_out_1192;
  (* register *) pwire FA_out_1193;
  (* register *) pwire FA_out_1194;
  (* register *) pwire FA_out_1195;
  (* register *) pwire FA_out_1196;
  (* register *) pwire FA_out_1197;
  (* register *) pwire FA_out_1198;
  (* register *) pwire FA_out_1199;
  (* register *) pwire FA_out_1200;
  (* register *) pwire FA_out_1201;
  (* register *) pwire FA_out_1202;
  (* register *) pwire FA_out_1203;
  (* register *) pwire FA_out_1204;
  (* register *) pwire FA_out_1205;
  (* register *) pwire FA_out_1206;
  (* register *) pwire FA_out_1207;
  (* register *) pwire FA_out_1208;
  (* register *) pwire FA_out_1209;
  (* register *) pwire FA_out_1210;
  (* register *) pwire FA_out_1211;
  (* register *) pwire FA_out_1212;
  (* register *) pwire FA_out_1213;
  (* register *) pwire FA_out_1214;
  (* register *) pwire FA_out_1215;
  (* register *) pwire FA_out_1216;
  (* register *) pwire FA_out_1217;
  (* register *) pwire FA_out_1218;
  (* register *) pwire FA_out_1219;
  (* register *) pwire FA_out_1220;
  (* register *) pwire FA_out_1221;
  (* register *) pwire FA_out_1222;
  (* register *) pwire FA_out_1223;
  (* register *) pwire FA_out_1224;
  (* register *) pwire FA_out_1225;
  (* register *) pwire FA_out_1226;
  (* register *) pwire FA_out_1227;
  (* register *) pwire FA_out_1228;
  (* register *) pwire FA_out_1229;
  (* register *) pwire FA_out_1230;
  (* register *) pwire FA_out_1231;
  (* register *) pwire FA_out_1232;
  (* register *) pwire FA_out_1233;
  (* register *) pwire FA_out_1234;
  (* register *) pwire FA_out_1235;
  (* register *) pwire FA_out_1236;
  (* register *) pwire FA_out_1237;
  (* register *) pwire FA_out_1238;
  (* register *) pwire FA_out_1239;
  (* register *) pwire FA_out_1240;
  (* register *) pwire FA_out_1241;
  (* register *) pwire FA_out_1242;
  (* register *) pwire FA_out_1243;
  (* register *) pwire FA_out_1244;
  (* register *) pwire FA_out_1245;
  (* register *) pwire FA_out_1246;
  (* register *) pwire FA_out_1247;
  (* register *) pwire FA_out_1248;
  (* register *) pwire FA_out_1249;
  (* register *) pwire FA_out_1250;
  (* register *) pwire FA_out_1251;
  (* register *) pwire FA_out_1252;
  (* register *) pwire FA_out_1253;
  (* register *) pwire FA_out_1254;
  (* register *) pwire FA_out_1255;
  (* register *) pwire FA_out_1256;
  (* register *) pwire FA_out_1257;
  (* register *) pwire FA_out_1258;
  (* register *) pwire FA_out_1259;
  (* register *) pwire FA_out_1260;
  (* register *) pwire FA_out_1261;
  (* register *) pwire FA_out_1262;
  (* register *) pwire FA_out_1263;
  (* register *) pwire FA_out_1264;
  (* register *) pwire FA_out_1265;
  (* register *) pwire FA_out_1266;
  (* register *) pwire FA_out_1267;
  (* register *) pwire FA_out_1268;
  (* register *) pwire FA_out_1269;
  (* register *) pwire FA_out_1270;
  (* register *) pwire FA_out_1271;
  (* register *) pwire FA_out_1272;
  (* register *) pwire FA_out_1273;
  (* register *) pwire FA_out_1274;
  (* register *) pwire FA_out_1275;
  (* register *) pwire FA_out_1276;
  (* register *) pwire FA_out_1277;
  (* register *) pwire FA_out_1278;
  (* register *) pwire FA_out_1279;
  (* register *) pwire FA_out_1280;
  (* register *) pwire FA_out_1281;
  (* register *) pwire FA_out_1282;
  (* register *) pwire FA_out_1283;
  (* register *) pwire FA_out_1284;
  (* register *) pwire FA_out_1285;
  (* register *) pwire FA_out_1286;
  (* register *) pwire FA_out_1287;
  (* register *) pwire FA_out_1288;
  (* register *) pwire FA_out_1289;
  (* register *) pwire FA_out_1290;
  (* register *) pwire FA_out_1291;
  (* register *) pwire FA_out_1292;
  (* register *) pwire FA_out_1293;
  (* register *) pwire FA_out_1294;
  (* register *) pwire FA_out_1295;
  (* register *) pwire FA_out_1296;
  (* register *) pwire FA_out_1297;
  (* register *) pwire FA_out_1298;
  (* register *) pwire FA_out_1299;
  (* register *) pwire FA_out_1300;
  (* register *) pwire FA_out_1301;
  (* register *) pwire FA_out_1302;
  (* register *) pwire FA_out_1303;
  (* register *) pwire FA_out_1304;
  (* register *) pwire FA_out_1305;
  (* register *) pwire FA_out_1306;
  (* register *) pwire FA_out_1307;
  (* register *) pwire FA_out_1308;
  (* register *) pwire FA_out_1309;
  (* register *) pwire FA_out_1310;
  (* register *) pwire FA_out_1311;
  (* register *) pwire FA_out_1312;
  (* register *) pwire FA_out_1313;
  (* register *) pwire FA_out_1314;
  (* register *) pwire FA_out_1315;
  (* register *) pwire FA_out_1316;
  (* register *) pwire FA_out_1317;
  (* register *) pwire FA_out_1318;
  (* register *) pwire FA_out_1319;
  (* register *) pwire FA_out_1320;
  (* register *) pwire FA_out_1321;
  (* register *) pwire FA_out_1322;
  (* register *) pwire FA_out_1323;
  (* register *) pwire FA_out_1324;
  (* register *) pwire FA_out_1325;
  (* register *) pwire FA_out_1326;
  (* register *) pwire FA_out_1327;
  (* register *) pwire FA_out_1328;
  (* register *) pwire FA_out_1329;
  (* register *) pwire FA_out_1330;
  (* register *) pwire FA_out_1331;
  (* register *) pwire FA_out_1332;
  (* register *) pwire FA_out_1333;
  (* register *) pwire FA_out_1334;
  (* register *) pwire FA_out_1335;
  (* register *) pwire FA_out_1336;
  (* register *) pwire FA_out_1337;
  (* register *) pwire FA_out_1338;
  (* register *) pwire FA_out_1339;
  (* register *) pwire FA_out_1340;
  (* register *) pwire FA_out_1341;
  (* register *) pwire FA_out_1342;
  (* register *) pwire FA_out_1343;
  (* register *) pwire FA_out_1344;
  (* register *) pwire FA_out_1345;
  (* register *) pwire FA_out_1346;
  (* register *) pwire FA_out_1347;
  (* register *) pwire FA_out_1348;
  (* register *) pwire FA_out_1349;
  (* register *) pwire FA_out_1350;
  (* register *) pwire FA_out_1351;
  (* register *) pwire FA_out_1352;
  (* register *) pwire FA_out_1353;
  (* register *) pwire FA_out_1354;
  (* register *) pwire FA_out_1355;
  (* register *) pwire FA_out_1356;
  (* register *) pwire FA_out_1357;
  (* register *) pwire FA_out_1358;
  (* register *) pwire FA_out_1359;
  (* register *) pwire FA_out_1360;
  (* register *) pwire FA_out_1361;
  (* register *) pwire FA_out_1362;
  (* register *) pwire FA_out_1363;
  (* register *) pwire FA_out_1364;
  (* register *) pwire FA_out_1365;
  (* register *) pwire FA_out_1366;
  (* register *) pwire FA_out_1367;
  (* register *) pwire FA_out_1368;
  (* register *) pwire FA_out_1369;
  (* register *) pwire FA_out_1370;
  (* register *) pwire FA_out_1371;
  (* register *) pwire FA_out_1372;
  (* register *) pwire FA_out_1373;
  (* register *) pwire FA_out_1374;
  (* register *) pwire FA_out_1375;
  (* register *) pwire FA_out_1376;
  (* register *) pwire FA_out_1377;
  (* register *) pwire FA_out_1378;
  (* register *) pwire FA_out_1379;
  (* register *) pwire FA_out_1380;
  (* register *) pwire FA_out_1381;
  (* register *) pwire FA_out_1382;
  (* register *) pwire FA_out_1383;
  (* register *) pwire FA_out_1384;
  (* register *) pwire FA_out_1385;
  (* register *) pwire FA_out_1386;
  (* register *) pwire FA_out_1387;
  (* register *) pwire FA_out_1388;
  (* register *) pwire FA_out_1389;
  (* register *) pwire FA_out_1390;
  (* register *) pwire FA_out_1391;
  (* register *) pwire FA_out_1392;
  (* register *) pwire FA_out_1393;
  (* register *) pwire FA_out_1394;
  (* register *) pwire FA_out_1395;
  (* register *) pwire FA_out_1396;
  (* register *) pwire FA_out_1397;
  (* register *) pwire FA_out_1398;
  (* register *) pwire FA_out_1399;
  (* register *) pwire FA_out_1400;
  (* register *) pwire FA_out_1401;
  (* register *) pwire FA_out_1402;
  (* register *) pwire FA_out_1403;
  (* register *) pwire FA_out_1404;
  (* register *) pwire FA_out_1405;
  (* register *) pwire FA_out_1406;
  (* register *) pwire FA_out_1407;
  (* register *) pwire FA_out_1408;
  (* register *) pwire FA_out_1409;
  (* register *) pwire FA_out_1410;
  (* register *) pwire FA_out_1411;
  (* register *) pwire FA_out_1412;
  (* register *) pwire FA_out_1413;
  (* register *) pwire FA_out_1414;
  (* register *) pwire FA_out_1415;
  (* register *) pwire FA_out_1416;
  (* register *) pwire FA_out_1417;
  (* register *) pwire FA_out_1418;
  (* register *) pwire FA_out_1419;
  (* register *) pwire FA_out_1420;
  (* register *) pwire FA_out_1421;
  (* register *) pwire FA_out_1422;
  (* register *) pwire FA_out_1423;
  (* register *) pwire FA_out_1424;
  (* register *) pwire FA_out_1425;
  (* register *) pwire FA_out_1426;
  (* register *) pwire FA_out_1427;
  (* register *) pwire FA_out_1428;
  (* register *) pwire FA_out_1429;
  (* register *) pwire FA_out_1430;
  (* register *) pwire FA_out_1431;
  (* register *) pwire FA_out_1432;
  (* register *) pwire FA_out_1433;
  (* register *) pwire FA_out_1434;
  (* register *) pwire FA_out_1435;
  (* register *) pwire FA_out_1436;
  (* register *) pwire FA_out_1437;
  (* register *) pwire FA_out_1438;
  (* register *) pwire FA_out_1439;
  (* register *) pwire FA_out_1440;
  (* register *) pwire FA_out_1441;
  (* register *) pwire FA_out_1442;
  (* register *) pwire FA_out_1443;
  (* register *) pwire FA_out_1444;
  (* register *) pwire FA_out_1445;
  (* register *) pwire FA_out_1446;
  (* register *) pwire FA_out_1447;
  (* register *) pwire FA_out_1448;
  (* register *) pwire FA_out_1449;
  (* register *) pwire FA_out_1450;
  (* register *) pwire FA_out_1451;
  (* register *) pwire FA_out_1452;
  (* register *) pwire FA_out_1453;
  (* register *) pwire FA_out_1454;
  (* register *) pwire FA_out_1455;
  (* register *) pwire FA_out_1456;
  (* register *) pwire FA_out_1457;
  (* register *) pwire FA_out_1458;
  (* register *) pwire FA_out_1459;
  (* register *) pwire FA_out_1460;
  (* register *) pwire FA_out_1461;
  (* register *) pwire FA_out_1462;
  (* register *) pwire FA_out_1463;
  (* register *) pwire FA_out_1464;
  (* register *) pwire FA_out_1465;
  (* register *) pwire FA_out_1466;
  (* register *) pwire FA_out_1467;
  (* register *) pwire FA_out_1468;
  (* register *) pwire FA_out_1469;
  (* register *) pwire FA_out_1470;
  (* register *) pwire FA_out_1471;
  (* register *) pwire FA_out_1472;
  (* register *) pwire FA_out_1473;
  (* register *) pwire FA_out_1474;
  (* register *) pwire FA_out_1475;
  (* register *) pwire FA_out_1476;
  (* register *) pwire FA_out_1477;
  (* register *) pwire FA_out_1478;
  (* register *) pwire FA_out_1479;
  (* register *) pwire FA_out_1480;
  (* register *) pwire FA_out_1481;
  (* register *) pwire FA_out_1482;
  (* register *) pwire FA_out_1483;
  (* register *) pwire FA_out_1484;
  (* register *) pwire FA_out_1485;
  (* register *) pwire FA_out_1486;
  (* register *) pwire FA_out_1487;
  (* register *) pwire FA_out_1488;
  (* register *) pwire FA_out_1489;
  (* register *) pwire FA_out_1490;
  (* register *) pwire FA_out_1491;
  (* register *) pwire FA_out_1492;
  (* register *) pwire FA_out_1493;
  (* register *) pwire FA_out_1494;
  (* register *) pwire FA_out_1495;
  (* register *) pwire FA_out_1496;
  (* register *) pwire FA_out_1497;
  (* register *) pwire FA_out_1498;
  (* register *) pwire FA_out_1499;
  (* register *) pwire FA_out_1500;
  (* register *) pwire FA_out_1501;
  (* register *) pwire FA_out_1502;
  (* register *) pwire FA_out_1503;
  (* register *) pwire FA_out_1504;
  (* register *) pwire FA_out_1505;
  (* register *) pwire FA_out_1506;
  (* register *) pwire FA_out_1507;
  (* register *) pwire FA_out_1508;
  (* register *) pwire FA_out_1509;
  (* register *) pwire FA_out_1510;
  (* register *) pwire FA_out_1511;
  (* register *) pwire FA_out_1512;
  (* register *) pwire FA_out_1513;
  (* register *) pwire FA_out_1514;
  (* register *) pwire FA_out_1515;
  (* register *) pwire FA_out_1516;
  (* register *) pwire FA_out_1517;
  (* register *) pwire FA_out_1518;
  (* register *) pwire FA_out_1519;
  (* register *) pwire FA_out_1520;
  (* register *) pwire FA_out_1521;
  (* register *) pwire FA_out_1522;
  (* register *) pwire FA_out_1523;
  (* register *) pwire FA_out_1524;
  (* register *) pwire FA_out_1525;
  (* register *) pwire FA_out_1526;
  (* register *) pwire FA_out_1527;
  (* register *) pwire FA_out_1528;
  (* register *) pwire FA_out_1529;
  (* register *) pwire FA_out_1530;
  (* register *) pwire FA_out_1531;
  (* register *) pwire FA_out_1532;
  (* register *) pwire FA_out_1533;
  (* register *) pwire FA_out_1534;
  (* register *) pwire FA_out_1535;
  (* register *) pwire FA_out_1536;
  (* register *) pwire FA_out_1537;
  (* register *) pwire FA_out_1538;
  (* register *) pwire FA_out_1539;
  (* register *) pwire FA_out_1540;
  (* register *) pwire FA_out_1541;
  (* register *) pwire FA_out_1542;
  (* register *) pwire FA_out_1543;
  (* register *) pwire FA_out_1544;
  (* register *) pwire FA_out_1545;
  (* register *) pwire FA_out_1546;
  (* register *) pwire FA_out_1547;
  (* register *) pwire FA_out_1548;
  (* register *) pwire FA_out_1549;
  (* register *) pwire FA_out_1550;
  (* register *) pwire FA_out_1551;
  (* register *) pwire FA_out_1552;
  (* register *) pwire FA_out_1553;
  (* register *) pwire FA_out_1554;
  (* register *) pwire FA_out_1555;
  (* register *) pwire FA_out_1556;
  (* register *) pwire FA_out_1557;
  (* register *) pwire FA_out_1558;
  (* register *) pwire FA_out_1559;
  (* register *) pwire FA_out_1560;
  (* register *) pwire FA_out_1561;
  (* register *) pwire FA_out_1562;
  (* register *) pwire FA_out_1563;
  (* register *) pwire FA_out_1564;
  (* register *) pwire FA_out_1565;
  (* register *) pwire FA_out_1566;
  (* register *) pwire FA_out_1567;
  (* register *) pwire FA_out_1568;
  (* register *) pwire FA_out_1569;
  (* register *) pwire FA_out_1570;
  (* register *) pwire FA_out_1571;
  (* register *) pwire FA_out_1572;
  (* register *) pwire FA_out_1573;
  (* register *) pwire FA_out_1574;
  (* register *) pwire FA_out_1575;
  (* register *) pwire FA_out_1576;
  (* register *) pwire FA_out_1577;
  (* register *) pwire FA_out_1578;
  (* register *) pwire FA_out_1579;
  (* register *) pwire FA_out_1580;
  (* register *) pwire FA_out_1581;
  (* register *) pwire FA_out_1582;
  (* register *) pwire FA_out_1583;
  (* register *) pwire FA_out_1584;
  (* register *) pwire FA_out_1585;
  (* register *) pwire FA_out_1586;
  (* register *) pwire FA_out_1587;
  (* register *) pwire FA_out_1588;
  (* register *) pwire FA_out_1589;
  (* register *) pwire FA_out_1590;
  (* register *) pwire FA_out_1591;
  (* register *) pwire FA_out_1592;
  (* register *) pwire FA_out_1593;
  (* register *) pwire FA_out_1594;
  (* register *) pwire FA_out_1595;
  (* register *) pwire FA_out_1596;
  (* register *) pwire FA_out_1597;
  (* register *) pwire FA_out_1598;
  (* register *) pwire FA_out_1599;
  (* register *) pwire FA_out_1600;
  (* register *) pwire FA_out_1601;
  (* register *) pwire FA_out_1602;
  (* register *) pwire FA_out_1603;
  (* register *) pwire FA_out_1604;
  (* register *) pwire FA_out_1605;
  (* register *) pwire FA_out_1606;
  (* register *) pwire FA_out_1607;
  (* register *) pwire FA_out_1608;
  (* register *) pwire FA_out_1609;
  (* register *) pwire FA_out_1610;
  (* register *) pwire FA_out_1611;
  (* register *) pwire FA_out_1612;
  (* register *) pwire FA_out_1613;
  (* register *) pwire FA_out_1614;
  (* register *) pwire FA_out_1615;
  (* register *) pwire FA_out_1616;
  (* register *) pwire FA_out_1617;
  (* register *) pwire FA_out_1618;
  (* register *) pwire FA_out_1619;
  (* register *) pwire FA_out_1620;
  (* register *) pwire FA_out_1621;
  (* register *) pwire FA_out_1622;
  (* register *) pwire FA_out_1623;
  (* register *) pwire FA_out_1624;
  (* register *) pwire FA_out_1625;
  (* register *) pwire FA_out_1626;
  (* register *) pwire FA_out_1627;
  (* register *) pwire FA_out_1628;
  (* register *) pwire FA_out_1629;
  (* register *) pwire FA_out_1630;
  (* register *) pwire FA_out_1631;
  (* register *) pwire FA_out_1632;
  (* register *) pwire FA_out_1633;
  (* register *) pwire FA_out_1634;
  (* register *) pwire FA_out_1635;
  (* register *) pwire FA_out_1636;
  (* register *) pwire FA_out_1637;
  (* register *) pwire FA_out_1638;
  (* register *) pwire FA_out_1639;
  (* register *) pwire FA_out_1640;
  (* register *) pwire FA_out_1641;
  (* register *) pwire FA_out_1642;
  (* register *) pwire FA_out_1643;
  (* register *) pwire FA_out_1644;
  (* register *) pwire FA_out_1645;
  (* register *) pwire FA_out_1646;
  (* register *) pwire FA_out_1647;
  (* register *) pwire FA_out_1648;
  (* register *) pwire FA_out_1649;
  (* register *) pwire FA_out_1650;
  (* register *) pwire FA_out_1651;
  (* register *) pwire FA_out_1652;
  (* register *) pwire FA_out_1653;
  (* register *) pwire FA_out_1654;
  (* register *) pwire FA_out_1655;
  (* register *) pwire FA_out_1656;
  (* register *) pwire FA_out_1657;
  (* register *) pwire FA_out_1658;
  (* register *) pwire FA_out_1659;
  (* register *) pwire FA_out_1660;
  (* register *) pwire FA_out_1661;
  (* register *) pwire FA_out_1662;
  (* register *) pwire FA_out_1663;
  (* register *) pwire FA_out_1664;
  (* register *) pwire FA_out_1665;
  (* register *) pwire FA_out_1666;
  (* register *) pwire FA_out_1667;
  (* register *) pwire FA_out_1668;
  (* register *) pwire FA_out_1669;
  (* register *) pwire FA_out_1670;
  (* register *) pwire FA_out_1671;
  (* register *) pwire FA_out_1672;
  (* register *) pwire FA_out_1673;
  (* register *) pwire FA_out_1674;
  (* register *) pwire FA_out_1675;
  (* register *) pwire FA_out_1676;
  (* register *) pwire FA_out_1677;
  (* register *) pwire FA_out_1678;
  (* register *) pwire FA_out_1679;
  (* register *) pwire FA_out_1680;
  (* register *) pwire FA_out_1681;
  (* register *) pwire FA_out_1682;
  (* register *) pwire FA_out_1683;
  (* register *) pwire FA_out_1684;
  (* register *) pwire FA_out_1685;
  (* register *) pwire FA_out_1686;
  (* register *) pwire FA_out_1687;
  (* register *) pwire FA_out_1688;
  (* register *) pwire FA_out_1689;
  (* register *) pwire FA_out_1690;
  (* register *) pwire FA_out_1691;
  (* register *) pwire FA_out_1692;
  (* register *) pwire FA_out_1693;
  (* register *) pwire FA_out_1694;
  (* register *) pwire FA_out_1695;
  (* register *) pwire FA_out_1696;
  (* register *) pwire FA_out_1697;
  (* register *) pwire FA_out_1698;
  (* register *) pwire FA_out_1699;
  (* register *) pwire FA_out_1700;
  (* register *) pwire FA_out_1701;
  (* register *) pwire FA_out_1702;
  (* register *) pwire FA_out_1703;
  (* register *) pwire FA_out_1704;
  (* register *) pwire FA_out_1705;
  (* register *) pwire FA_out_1706;
  (* register *) pwire FA_out_1707;
  (* register *) pwire FA_out_1708;
  (* register *) pwire FA_out_1709;
  (* register *) pwire FA_out_1710;
  (* register *) pwire FA_out_1711;
  (* register *) pwire FA_out_1712;
  (* register *) pwire FA_out_1713;
  (* register *) pwire FA_out_1714;
  (* register *) pwire FA_out_1715;
  (* register *) pwire FA_out_1716;
  (* register *) pwire FA_out_1717;
  (* register *) pwire FA_out_1718;
  (* register *) pwire FA_out_1719;
  (* register *) pwire FA_out_1720;
  (* register *) pwire FA_out_1721;
  (* register *) pwire FA_out_1722;
  (* register *) pwire FA_out_1723;
  (* register *) pwire FA_out_1724;
  (* register *) pwire FA_out_1725;
  (* register *) pwire FA_out_1726;
  (* register *) pwire FA_out_1727;
  (* register *) pwire FA_out_1728;
  (* register *) pwire FA_out_1729;
  (* register *) pwire FA_out_1730;
  (* register *) pwire FA_out_1731;
  (* register *) pwire FA_out_1732;
  (* register *) pwire FA_out_1733;
  (* register *) pwire FA_out_1734;
  (* register *) pwire FA_out_1735;
  (* register *) pwire FA_out_1736;
  (* register *) pwire FA_out_1737;
  (* register *) pwire FA_out_1738;
  (* register *) pwire FA_out_1739;
  (* register *) pwire FA_out_1740;
  (* register *) pwire FA_out_1741;
  (* register *) pwire FA_out_1742;
  (* register *) pwire FA_out_1743;
  (* register *) pwire FA_out_1744;
  (* register *) pwire FA_out_1745;
  (* register *) pwire FA_out_1746;
  (* register *) pwire FA_out_1747;
  (* register *) pwire FA_out_1748;
  (* register *) pwire FA_out_1749;
  (* register *) pwire FA_out_1750;
  (* register *) pwire FA_out_1751;
  (* register *) pwire FA_out_1752;
  (* register *) pwire FA_out_1753;
  (* register *) pwire FA_out_1754;
  (* register *) pwire FA_out_1755;
  (* register *) pwire FA_out_1756;
  (* register *) pwire FA_out_1757;
  (* register *) pwire FA_out_1758;
  (* register *) pwire FA_out_1759;
  (* register *) pwire FA_out_1760;
  (* register *) pwire FA_out_1761;
  (* register *) pwire FA_out_1762;
  (* register *) pwire FA_out_1763;
  (* register *) pwire FA_out_1764;
  (* register *) pwire FA_out_1765;
  (* register *) pwire FA_out_1766;
  (* register *) pwire FA_out_1767;
  (* register *) pwire FA_out_1768;
  (* register *) pwire FA_out_1769;
  (* register *) pwire FA_out_1770;
  (* register *) pwire FA_out_1771;
  (* register *) pwire FA_out_1772;
  (* register *) pwire FA_out_1773;
  (* register *) pwire FA_out_1774;
  (* register *) pwire FA_out_1775;
  (* register *) pwire FA_out_1776;
  (* register *) pwire FA_out_1777;
  (* register *) pwire FA_out_1778;
  (* register *) pwire FA_out_1779;
  (* register *) pwire FA_out_1780;
  (* register *) pwire FA_out_1781;
  (* register *) pwire FA_out_1782;
  (* register *) pwire FA_out_1783;
  (* register *) pwire FA_out_1784;
  (* register *) pwire FA_out_1785;
  (* register *) pwire FA_out_1786;
  (* register *) pwire FA_out_1787;
  (* register *) pwire FA_out_1788;
  (* register *) pwire FA_out_1789;
  (* register *) pwire FA_out_1790;
  (* register *) pwire FA_out_1791;
  (* register *) pwire FA_out_1792;
  (* register *) pwire FA_out_1793;
  (* register *) pwire FA_out_1794;
  (* register *) pwire FA_out_1795;
  (* register *) pwire FA_out_1796;
  (* register *) pwire FA_out_1797;
  (* register *) pwire FA_out_1798;
  (* register *) pwire FA_out_1799;
  (* register *) pwire FA_out_1800;
  (* register *) pwire FA_out_1801;
  (* register *) pwire FA_out_1802;
  (* register *) pwire FA_out_1803;
  (* register *) pwire FA_out_1804;
  (* register *) pwire FA_out_1805;
  (* register *) pwire FA_out_1806;
  (* register *) pwire FA_out_1807;
  (* register *) pwire FA_out_1808;
  (* register *) pwire FA_out_1809;
  (* register *) pwire FA_out_1810;
  (* register *) pwire FA_out_1811;
  (* register *) pwire FA_out_1812;
  (* register *) pwire FA_out_1813;
  (* register *) pwire FA_out_1814;
  (* register *) pwire FA_out_1815;
  (* register *) pwire FA_out_1816;
  (* register *) pwire FA_out_1817;
  (* register *) pwire FA_out_1818;
  (* register *) pwire FA_out_1819;
  (* register *) pwire FA_out_1820;
  (* register *) pwire FA_out_1821;
  (* register *) pwire FA_out_1822;
  (* register *) pwire FA_out_1823;
  (* register *) pwire FA_out_1824;
  (* register *) pwire FA_out_1825;
  (* register *) pwire FA_out_1826;
  (* register *) pwire FA_out_1827;
  (* register *) pwire FA_out_1828;
  (* register *) pwire FA_out_1829;
  (* register *) pwire FA_out_1830;
  (* register *) pwire FA_out_1831;
  (* register *) pwire FA_out_1832;
  (* register *) pwire FA_out_1833;
  (* register *) pwire FA_out_1834;
  (* register *) pwire FA_out_1835;
  (* register *) pwire FA_out_1836;
  (* register *) pwire FA_out_1837;
  (* register *) pwire FA_out_1838;
  (* register *) pwire FA_out_1839;
  (* register *) pwire FA_out_1840;
  (* register *) pwire FA_out_1841;
  (* register *) pwire FA_out_1842;
  (* register *) pwire FA_out_1843;
  (* register *) pwire FA_out_1844;
  (* register *) pwire FA_out_1845;
  (* register *) pwire FA_out_1846;
  (* register *) pwire FA_out_1847;
  (* register *) pwire FA_out_1848;
  (* register *) pwire FA_out_1849;
  (* register *) pwire FA_out_1850;
  (* register *) pwire FA_out_1851;
  (* register *) pwire FA_out_1852;
  (* register *) pwire FA_out_1853;
  (* register *) pwire FA_out_1854;
  (* register *) pwire FA_out_1855;
  (* register *) pwire FA_out_1856;
  (* register *) pwire FA_out_1857;
  (* register *) pwire FA_out_1858;
  (* register *) pwire FA_out_1859;
  (* register *) pwire FA_out_1860;
  (* register *) pwire FA_out_1861;
  (* register *) pwire FA_out_1862;
  (* register *) pwire FA_out_1863;
  (* register *) pwire FA_out_1864;
  (* register *) pwire FA_out_1865;
  (* register *) pwire FA_out_1866;
  (* register *) pwire FA_out_1867;
  (* register *) pwire FA_out_1868;
  (* register *) pwire FA_out_1869;
  (* register *) pwire FA_out_1870;
  (* register *) pwire FA_out_1871;
  (* register *) pwire FA_out_1872;
  (* register *) pwire FA_out_1873;
  (* register *) pwire FA_out_1874;
  (* register *) pwire FA_out_1875;
  (* register *) pwire FA_out_1876;
  (* register *) pwire FA_out_1877;
  (* register *) pwire FA_out_1878;
  (* register *) pwire FA_out_1879;
  (* register *) pwire FA_out_1880;
  (* register *) pwire FA_out_1881;
  (* register *) pwire FA_out_1882;
  (* register *) pwire FA_out_1883;
  (* register *) pwire FA_out_1884;
  (* register *) pwire FA_out_1885;
  (* register *) pwire FA_out_1886;
  (* register *) pwire FA_out_1887;
  (* register *) pwire FA_out_1888;
  (* register *) pwire FA_out_1889;
  (* register *) pwire FA_out_1890;
  (* register *) pwire FA_out_1891;
  (* register *) pwire FA_out_1892;
  (* register *) pwire FA_out_1893;
  (* register *) pwire FA_out_1894;
  (* register *) pwire FA_out_1895;
  (* register *) pwire FA_out_1896;
  (* register *) pwire FA_out_1897;
  (* register *) pwire FA_out_1898;
  (* register *) pwire FA_out_1899;
  (* register *) pwire FA_out_1900;
  (* register *) pwire FA_out_1901;
  (* register *) pwire FA_out_1902;
  (* register *) pwire FA_out_1903;
  (* register *) pwire FA_out_1904;
  (* register *) pwire FA_out_1905;
  (* register *) pwire FA_out_1906;
  (* register *) pwire FA_out_1907;
  (* register *) pwire FA_out_1908;
  (* register *) pwire FA_out_1909;
  (* register *) pwire FA_out_1910;
  (* register *) pwire FA_out_1911;
  (* register *) pwire FA_out_1912;
  (* register *) pwire FA_out_1913;
  (* register *) pwire FA_out_1914;
  (* register *) pwire FA_out_1915;
  (* register *) pwire FA_out_1916;
  (* register *) pwire FA_out_1917;
  (* register *) pwire FA_out_1918;
  (* register *) pwire FA_out_1919;
  (* register *) pwire FA_out_1920;
  (* register *) pwire FA_out_1921;
  (* register *) pwire FA_out_1922;
  (* register *) pwire FA_out_1923;
  (* register *) pwire FA_out_1924;
  (* register *) pwire FA_out_1925;
  (* register *) pwire FA_out_1926;
  (* register *) pwire FA_out_1927;
  (* register *) pwire FA_out_1928;
  (* register *) pwire FA_out_1929;
  (* register *) pwire FA_out_1930;
  (* register *) pwire FA_out_1931;
  (* register *) pwire FA_out_1932;
  (* register *) pwire FA_out_1933;
  (* register *) pwire FA_out_1934;
  (* register *) pwire FA_out_1935;
  (* register *) pwire FA_out_1936;
  (* register *) pwire FA_out_1937;
  (* register *) pwire FA_out_1938;
  (* register *) pwire FA_out_1939;
  (* register *) pwire FA_out_1940;
  (* register *) pwire FA_out_1941;
  (* register *) pwire FA_out_1942;
  (* register *) pwire FA_out_1943;
  (* register *) pwire FA_out_1944;
  (* register *) pwire FA_out_1945;
  (* register *) pwire FA_out_1946;
  (* register *) pwire FA_out_1947;
  (* register *) pwire FA_out_1948;
  (* register *) pwire FA_out_1949;
  (* register *) pwire FA_out_1950;
  (* register *) pwire FA_out_1951;
  (* register *) pwire FA_out_1952;
  (* register *) pwire FA_out_1953;
  (* register *) pwire FA_out_1954;
  (* register *) pwire FA_out_1955;
  (* register *) pwire FA_out_1956;
  (* register *) pwire FA_out_1957;
  (* register *) pwire FA_out_1958;
  (* register *) pwire FA_out_1959;
  (* register *) pwire FA_out_1960;
  (* register *) pwire FA_out_1961;
  (* register *) pwire FA_out_1962;
  (* register *) pwire FA_out_1963;
  (* register *) pwire FA_out_1964;
  (* register *) pwire FA_out_1965;
  (* register *) pwire FA_out_1966;
  (* register *) pwire FA_out_1967;
  (* register *) pwire FA_out_1968;
  (* register *) pwire FA_out_1969;
  (* register *) pwire FA_out_1970;
  (* register *) pwire FA_out_1971;
  (* register *) pwire FA_out_1972;
  (* register *) pwire FA_out_1973;
  (* register *) pwire FA_out_1974;
  (* register *) pwire FA_out_1975;
  (* register *) pwire FA_out_1976;
  (* register *) pwire FA_out_1977;
  (* register *) pwire FA_out_1978;
  (* register *) pwire FA_out_1979;
  (* register *) pwire FA_out_1980;
  (* register *) pwire FA_out_1981;
  (* register *) pwire FA_out_1982;
  (* register *) pwire FA_out_1983;
  (* register *) pwire FA_out_1984;
  (* register *) pwire FA_out_1985;
  (* register *) pwire FA_out_1986;
  (* register *) pwire FA_out_1987;
  (* register *) pwire FA_out_1988;
  (* register *) pwire FA_out_1989;
  (* register *) pwire FA_out_1990;
  (* register *) pwire FA_out_1991;
  (* register *) pwire FA_out_1992;
  (* register *) pwire FA_out_1993;
  (* register *) pwire FA_out_1994;
  (* register *) pwire FA_out_1995;
  (* register *) pwire FA_out_1996;
  (* register *) pwire FA_out_1997;
  (* register *) pwire FA_out_1998;
  (* register *) pwire FA_out_1999;
  (* register *) pwire FA_out_2000;
  (* register *) pwire FA_out_2001;
  (* register *) pwire FA_out_2002;
  (* register *) pwire FA_out_2003;
  (* register *) pwire FA_out_2004;
  (* register *) pwire FA_out_2005;
  (* register *) pwire FA_out_2006;
  (* register *) pwire FA_out_2007;
  (* register *) pwire FA_out_2008;
  (* register *) pwire FA_out_2009;
  (* register *) pwire FA_out_2010;
  (* register *) pwire FA_out_2011;
  (* register *) pwire FA_out_2012;
  (* register *) pwire FA_out_2013;
  (* register *) pwire FA_out_2014;
  (* register *) pwire FA_out_2015;
  (* register *) pwire FA_out_2016;
  (* register *) pwire FA_out_2017;
  (* register *) pwire FA_out_2018;
  (* register *) pwire FA_out_2019;
  (* register *) pwire FA_out_2020;
  (* register *) pwire FA_out_2021;
  (* register *) pwire FA_out_2022;
  (* register *) pwire FA_out_2023;
  (* register *) pwire FA_out_2024;
  (* register *) pwire FA_out_2025;
  (* register *) pwire FA_out_2026;
  (* register *) pwire FA_out_2027;
  (* register *) pwire FA_out_2028;
  (* register *) pwire FA_out_2029;
  (* register *) pwire FA_out_2030;
  (* register *) pwire FA_out_2031;
  (* register *) pwire FA_out_2032;
  (* register *) pwire FA_out_2033;
  (* register *) pwire FA_out_2034;
  (* register *) pwire FA_out_2035;
  (* register *) pwire FA_out_2036;
  (* register *) pwire FA_out_2037;
  (* register *) pwire FA_out_2038;
  (* register *) pwire FA_out_2039;
  (* register *) pwire FA_out_2040;
  (* register *) pwire FA_out_2041;
  (* register *) pwire FA_out_2042;
  (* register *) pwire FA_out_2043;
  (* register *) pwire FA_out_2044;
  (* register *) pwire FA_out_2045;
  (* register *) pwire FA_out_2046;
  (* register *) pwire FA_out_2047;
  (* register *) pwire FA_out_2048;
  (* register *) pwire FA_out_2049;
  (* register *) pwire FA_out_2050;
  (* register *) pwire FA_out_2051;
  (* register *) pwire FA_out_2052;
  (* register *) pwire FA_out_2053;
  (* register *) pwire FA_out_2054;
  (* register *) pwire FA_out_2055;
  (* register *) pwire FA_out_2056;
  (* register *) pwire FA_out_2057;
  (* register *) pwire FA_out_2058;
  (* register *) pwire FA_out_2059;
  (* register *) pwire FA_out_2060;
  (* register *) pwire FA_out_2061;
  (* register *) pwire FA_out_2062;
  (* register *) pwire FA_out_2063;
  (* register *) pwire FA_out_2064;
  (* register *) pwire FA_out_2065;
  (* register *) pwire FA_out_2066;
  (* register *) pwire FA_out_2067;
  (* register *) pwire FA_out_2068;
  (* register *) pwire FA_out_2069;
  (* register *) pwire FA_out_2070;
  (* register *) pwire FA_out_2071;
  (* register *) pwire FA_out_2072;
  (* register *) pwire FA_out_2073;
  (* register *) pwire FA_out_2074;
  (* register *) pwire FA_out_2075;
  (* register *) pwire FA_out_2076;
  (* register *) pwire FA_out_2077;
  (* register *) pwire FA_out_2078;
  (* register *) pwire FA_out_2079;
  (* register *) pwire FA_out_2080;
  (* register *) pwire FA_out_2081;
  (* register *) pwire FA_out_2082;
  (* register *) pwire FA_out_2083;
  (* register *) pwire FA_out_2084;
  (* register *) pwire FA_out_2085;
  (* register *) pwire FA_out_2086;
  (* register *) pwire FA_out_2087;
  (* register *) pwire FA_out_2088;
  (* register *) pwire FA_out_2089;
  (* register *) pwire FA_out_2090;
  (* register *) pwire FA_out_2091;
  (* register *) pwire FA_out_2092;
  (* register *) pwire FA_out_2093;
  (* register *) pwire FA_out_2094;
  (* register *) pwire FA_out_2095;
  (* register *) pwire FA_out_2096;
  (* register *) pwire FA_out_2097;
  (* register *) pwire FA_out_2098;
  (* register *) pwire FA_out_2099;
  (* register *) pwire FA_out_2100;
  (* register *) pwire FA_out_2101;
  (* register *) pwire FA_out_2102;
  (* register *) pwire FA_out_2103;
  (* register *) pwire FA_out_2104;
  (* register *) pwire FA_out_2105;
  (* register *) pwire FA_out_2106;
  (* register *) pwire FA_out_2107;
  (* register *) pwire FA_out_2108;
  (* register *) pwire FA_out_2109;
  (* register *) pwire FA_out_2110;
  (* register *) pwire FA_out_2111;
  (* register *) pwire FA_out_2112;
  (* register *) pwire FA_out_2113;
  (* register *) pwire FA_out_2114;
  (* register *) pwire FA_out_2115;
  (* register *) pwire FA_out_2116;
  (* register *) pwire FA_out_2117;
  (* register *) pwire FA_out_2118;
  (* register *) pwire FA_out_2119;
  (* register *) pwire FA_out_2120;
  (* register *) pwire FA_out_2121;
  (* register *) pwire FA_out_2122;
  (* register *) pwire FA_out_2123;
  (* register *) pwire FA_out_2124;
  (* register *) pwire FA_out_2125;
  (* register *) pwire FA_out_2126;
  (* register *) pwire FA_out_2127;
  (* register *) pwire FA_out_2128;
  (* register *) pwire FA_out_2129;
  (* register *) pwire FA_out_2130;
  (* register *) pwire FA_out_2131;
  (* register *) pwire FA_out_2132;
  (* register *) pwire FA_out_2133;
  (* register *) pwire FA_out_2134;
  (* register *) pwire FA_out_2135;
  (* register *) pwire FA_out_2136;
  (* register *) pwire FA_out_2137;
  (* register *) pwire FA_out_2138;
  (* register *) pwire FA_out_2139;
  (* register *) pwire FA_out_2140;
  (* register *) pwire FA_out_2141;
  (* register *) pwire FA_out_2142;
  (* register *) pwire FA_out_2143;
  (* register *) pwire FA_out_2144;
  (* register *) pwire FA_out_2145;
  (* register *) pwire FA_out_2146;
  (* register *) pwire FA_out_2147;
  (* register *) pwire FA_out_2148;
  (* register *) pwire FA_out_2149;
  (* register *) pwire FA_out_2150;
  (* register *) pwire FA_out_2151;
  (* register *) pwire FA_out_2152;
  (* register *) pwire FA_out_2153;
  (* register *) pwire FA_out_2154;
  (* register *) pwire FA_out_2155;
  (* register *) pwire FA_out_2156;
  (* register *) pwire FA_out_2157;
  (* register *) pwire FA_out_2158;
  (* register *) pwire FA_out_2159;
  (* register *) pwire FA_out_2160;
  (* register *) pwire FA_out_2161;
  (* register *) pwire FA_out_2162;
  (* register *) pwire FA_out_2163;
  (* register *) pwire FA_out_2164;
  (* register *) pwire FA_out_2165;
  (* register *) pwire FA_out_2166;
  (* register *) pwire FA_out_2167;
  (* register *) pwire FA_out_2168;
  (* register *) pwire FA_out_2169;
  (* register *) pwire FA_out_2170;
  (* register *) pwire FA_out_2171;
  (* register *) pwire FA_out_2172;
  (* register *) pwire FA_out_2173;
  (* register *) pwire FA_out_2174;
  (* register *) pwire FA_out_2175;
  (* register *) pwire FA_out_2176;
  (* register *) pwire FA_out_2177;
  (* register *) pwire FA_out_2178;
  (* register *) pwire FA_out_2179;
  (* register *) pwire FA_out_2180;
  (* register *) pwire FA_out_2181;
  (* register *) pwire FA_out_2182;
  (* register *) pwire FA_out_2183;
  (* register *) pwire FA_out_2184;
  (* register *) pwire FA_out_2185;
  (* register *) pwire FA_out_2186;
  (* register *) pwire FA_out_2187;
  (* register *) pwire FA_out_2188;
  (* register *) pwire FA_out_2189;
  (* register *) pwire FA_out_2190;
  (* register *) pwire FA_out_2191;
  (* register *) pwire FA_out_2192;
  (* register *) pwire FA_out_2193;
  (* register *) pwire FA_out_2194;
  (* register *) pwire FA_out_2195;
  (* register *) pwire FA_out_2196;
  (* register *) pwire FA_out_2197;
  (* register *) pwire FA_out_2198;
  (* register *) pwire FA_out_2199;
  (* register *) pwire FA_out_2200;
  (* register *) pwire FA_out_2201;
  (* register *) pwire FA_out_2202;
  (* register *) pwire FA_out_2203;
  (* register *) pwire FA_out_2204;
  (* register *) pwire FA_out_2205;
  (* register *) pwire FA_out_2206;
  (* register *) pwire FA_out_2207;
  (* register *) pwire FA_out_2208;
  (* register *) pwire FA_out_2209;
  (* register *) pwire FA_out_2210;
  (* register *) pwire FA_out_2211;
  (* register *) pwire FA_out_2212;
  (* register *) pwire FA_out_2213;
  (* register *) pwire FA_out_2214;
  (* register *) pwire FA_out_2215;
  (* register *) pwire FA_out_2216;
  (* register *) pwire FA_out_2217;
  (* register *) pwire FA_out_2218;
  (* register *) pwire FA_out_2219;
  (* register *) pwire FA_out_2220;
  (* register *) pwire FA_out_2221;
  (* register *) pwire FA_out_2222;
  (* register *) pwire FA_out_2223;
  (* register *) pwire FA_out_2224;
  (* register *) pwire FA_out_2225;
  (* register *) pwire FA_out_2226;
  (* register *) pwire FA_out_2227;
  (* register *) pwire FA_out_2228;
  (* register *) pwire FA_out_2229;
  (* register *) pwire FA_out_2230;
  (* register *) pwire FA_out_2231;
  (* register *) pwire FA_out_2232;
  (* register *) pwire FA_out_2233;
  (* register *) pwire FA_out_2234;
  (* register *) pwire FA_out_2235;
  (* register *) pwire FA_out_2236;
  (* register *) pwire FA_out_2237;
  (* register *) pwire FA_out_2238;
  (* register *) pwire FA_out_2239;
  (* register *) pwire FA_out_2240;
  (* register *) pwire FA_out_2241;
  (* register *) pwire FA_out_2242;
  (* register *) pwire FA_out_2243;
  (* register *) pwire FA_out_2244;
  (* register *) pwire FA_out_2245;
  (* register *) pwire FA_out_2246;
  (* register *) pwire FA_out_2247;
  (* register *) pwire FA_out_2248;
  (* register *) pwire FA_out_2249;
  (* register *) pwire FA_out_2250;
  (* register *) pwire FA_out_2251;
  (* register *) pwire FA_out_2252;
  (* register *) pwire FA_out_2253;
  (* register *) pwire FA_out_2254;
  (* register *) pwire FA_out_2255;
  (* register *) pwire FA_out_2256;
  (* register *) pwire FA_out_2257;
  (* register *) pwire FA_out_2258;
  (* register *) pwire FA_out_2259;
  (* register *) pwire FA_out_2260;
  (* register *) pwire FA_out_2261;
  (* register *) pwire FA_out_2262;
  (* register *) pwire FA_out_2263;
  (* register *) pwire FA_out_2264;
  (* register *) pwire FA_out_2265;
  (* register *) pwire FA_out_2266;
  (* register *) pwire FA_out_2267;
  (* register *) pwire FA_out_2268;
  (* register *) pwire FA_out_2269;
  (* register *) pwire FA_out_2270;
  (* register *) pwire FA_out_2271;
  (* register *) pwire FA_out_2272;
  (* register *) pwire FA_out_2273;
  (* register *) pwire FA_out_2274;
  (* register *) pwire FA_out_2275;
  (* register *) pwire FA_out_2276;
  (* register *) pwire FA_out_2277;
  (* register *) pwire FA_out_2278;
  (* register *) pwire FA_out_2279;
  (* register *) pwire FA_out_2280;
  (* register *) pwire FA_out_2281;
  (* register *) pwire FA_out_2282;
  (* register *) pwire FA_out_2283;
  (* register *) pwire FA_out_2284;
  (* register *) pwire FA_out_2285;
  (* register *) pwire FA_out_2286;
  (* register *) pwire FA_out_2287;
  (* register *) pwire FA_out_2288;
  (* register *) pwire FA_out_2289;
  (* register *) pwire FA_out_2290;
  (* register *) pwire FA_out_2291;
  (* register *) pwire FA_out_2292;
  (* register *) pwire FA_out_2293;
  (* register *) pwire FA_out_2294;
  (* register *) pwire FA_out_2295;
  (* register *) pwire FA_out_2296;
  (* register *) pwire FA_out_2297;
  (* register *) pwire FA_out_2298;
  (* register *) pwire FA_out_2299;
  (* register *) pwire FA_out_2300;
  (* register *) pwire FA_out_2301;
  (* register *) pwire FA_out_2302;
  (* register *) pwire FA_out_2303;
  (* register *) pwire FA_out_2304;
  (* register *) pwire FA_out_2305;
  (* register *) pwire FA_out_2306;
  (* register *) pwire FA_out_2307;
  (* register *) pwire FA_out_2308;
  (* register *) pwire FA_out_2309;
  (* register *) pwire FA_out_2310;
  (* register *) pwire FA_out_2311;
  (* register *) pwire FA_out_2312;
  (* register *) pwire FA_out_2313;
  (* register *) pwire FA_out_2314;
  (* register *) pwire FA_out_2315;
  (* register *) pwire FA_out_2316;
  (* register *) pwire FA_out_2317;
  (* register *) pwire FA_out_2318;
  (* register *) pwire FA_out_2319;
  (* register *) pwire FA_out_2320;
  (* register *) pwire FA_out_2321;
  (* register *) pwire FA_out_2322;
  (* register *) pwire FA_out_2323;
  (* register *) pwire FA_out_2324;
  (* register *) pwire FA_out_2325;
  (* register *) pwire FA_out_2326;
  (* register *) pwire FA_out_2327;
  (* register *) pwire FA_out_2328;
  (* register *) pwire FA_out_2329;
  (* register *) pwire FA_out_2330;
  (* register *) pwire FA_out_2331;
  (* register *) pwire FA_out_2332;
  (* register *) pwire FA_out_2333;
  (* register *) pwire FA_out_2334;
  (* register *) pwire FA_out_2335;
  (* register *) pwire FA_out_2336;
  (* register *) pwire FA_out_2337;
  (* register *) pwire FA_out_2338;
  (* register *) pwire FA_out_2339;
  (* register *) pwire FA_out_2340;
  (* register *) pwire FA_out_2341;
  (* register *) pwire FA_out_2342;
  (* register *) pwire FA_out_2343;
  (* register *) pwire FA_out_2344;
  (* register *) pwire FA_out_2345;
  (* register *) pwire FA_out_2346;
  (* register *) pwire FA_out_2347;
  (* register *) pwire FA_out_2348;
  (* register *) pwire FA_out_2349;
  (* register *) pwire FA_out_2350;
  (* register *) pwire FA_out_2351;
  (* register *) pwire FA_out_2352;
  (* register *) pwire FA_out_2353;
  (* register *) pwire FA_out_2354;
  (* register *) pwire FA_out_2355;
  (* register *) pwire FA_out_2356;
  (* register *) pwire FA_out_2357;
  (* register *) pwire FA_out_2358;
  (* register *) pwire FA_out_2359;
  (* register *) pwire FA_out_2360;
  (* register *) pwire FA_out_2361;
  (* register *) pwire FA_out_2362;
  (* register *) pwire FA_out_2363;
  (* register *) pwire FA_out_2364;
  (* register *) pwire FA_out_2365;
  (* register *) pwire FA_out_2366;
  (* register *) pwire FA_out_2367;
  (* register *) pwire FA_out_2368;
  (* register *) pwire FA_out_2369;
  (* register *) pwire FA_out_2370;
  (* register *) pwire FA_out_2371;
  (* register *) pwire FA_out_2372;
  (* register *) pwire FA_out_2373;
  (* register *) pwire FA_out_2374;
  (* register *) pwire FA_out_2375;
  (* register *) pwire FA_out_2376;
  (* register *) pwire FA_out_2377;
  (* register *) pwire FA_out_2378;
  (* register *) pwire FA_out_2379;
  (* register *) pwire FA_out_2380;
  (* register *) pwire FA_out_2381;
  (* register *) pwire FA_out_2382;
  (* register *) pwire FA_out_2383;
  (* register *) pwire FA_out_2384;
  (* register *) pwire FA_out_2385;
  (* register *) pwire FA_out_2386;
  (* register *) pwire FA_out_2387;
  (* register *) pwire FA_out_2388;
  (* register *) pwire FA_out_2389;
  (* register *) pwire FA_out_2390;
  (* register *) pwire FA_out_2391;
  (* register *) pwire FA_out_2392;
  (* register *) pwire FA_out_2393;
  (* register *) pwire FA_out_2394;
  (* register *) pwire FA_out_2395;
  (* register *) pwire FA_out_2396;
  (* register *) pwire FA_out_2397;
  (* register *) pwire FA_out_2398;
  (* register *) pwire FA_out_2399;
  (* register *) pwire FA_out_2400;
  (* register *) pwire FA_out_2401;
  (* register *) pwire FA_out_2402;
  (* register *) pwire FA_out_2403;
  (* register *) pwire FA_out_2404;
  (* register *) pwire FA_out_2405;
  (* register *) pwire FA_out_2406;
  (* register *) pwire FA_out_2407;
  (* register *) pwire FA_out_2408;
  (* register *) pwire FA_out_2409;
  (* register *) pwire FA_out_2410;
  (* register *) pwire FA_out_2411;
  (* register *) pwire FA_out_2412;
  (* register *) pwire FA_out_2413;
  (* register *) pwire FA_out_2414;
  (* register *) pwire FA_out_2415;
  (* register *) pwire FA_out_2416;
  (* register *) pwire FA_out_2417;
  (* register *) pwire FA_out_2418;
  (* register *) pwire FA_out_2419;
  (* register *) pwire FA_out_2420;
  (* register *) pwire FA_out_2421;
  (* register *) pwire FA_out_2422;
  (* register *) pwire FA_out_2423;
  (* register *) pwire FA_out_2424;
  (* register *) pwire FA_out_2425;
  (* register *) pwire FA_out_2426;
  (* register *) pwire FA_out_2427;
  (* register *) pwire FA_out_2428;
  (* register *) pwire FA_out_2429;
  (* register *) pwire FA_out_2430;
  (* register *) pwire FA_out_2431;
  (* register *) pwire FA_out_2432;
  (* register *) pwire FA_out_2433;
  (* register *) pwire FA_out_2434;
  (* register *) pwire FA_out_2435;
  (* register *) pwire FA_out_2436;
  (* register *) pwire FA_out_2437;
  (* register *) pwire FA_out_2438;
  (* register *) pwire FA_out_2439;
  (* register *) pwire FA_out_2440;
  (* register *) pwire FA_out_2441;
  (* register *) pwire FA_out_2442;
  (* register *) pwire FA_out_2443;
  (* register *) pwire FA_out_2444;
  (* register *) pwire FA_out_2445;
  (* register *) pwire FA_out_2446;
  (* register *) pwire FA_out_2447;
  (* register *) pwire FA_out_2448;
  (* register *) pwire FA_out_2449;
  (* register *) pwire FA_out_2450;
  (* register *) pwire FA_out_2451;
  (* register *) pwire FA_out_2452;
  (* register *) pwire FA_out_2453;
  (* register *) pwire FA_out_2454;
  (* register *) pwire FA_out_2455;
  (* register *) pwire FA_out_2456;
  (* register *) pwire FA_out_2457;
  (* register *) pwire FA_out_2458;
  (* register *) pwire FA_out_2459;
  (* register *) pwire FA_out_2460;
  (* register *) pwire FA_out_2461;
  (* register *) pwire FA_out_2462;
  (* register *) pwire FA_out_2463;
  (* register *) pwire FA_out_2464;
  (* register *) pwire FA_out_2465;
  (* register *) pwire FA_out_2466;
  (* register *) pwire FA_out_2467;
  (* register *) pwire FA_out_2468;
  (* register *) pwire FA_out_2469;
  (* register *) pwire FA_out_2470;
  (* register *) pwire FA_out_2471;
  (* register *) pwire FA_out_2472;
  (* register *) pwire FA_out_2473;
  (* register *) pwire FA_out_2474;
  (* register *) pwire FA_out_2475;
  (* register *) pwire FA_out_2476;
  (* register *) pwire FA_out_2477;
  (* register *) pwire FA_out_2478;
  (* register *) pwire FA_out_2479;
  (* register *) pwire FA_out_2480;
  (* register *) pwire FA_out_2481;
  (* register *) pwire FA_out_2482;
  (* register *) pwire FA_out_2483;
  (* register *) pwire FA_out_2484;
  (* register *) pwire FA_out_2485;
  (* register *) pwire FA_out_2486;
  (* register *) pwire FA_out_2487;
  (* register *) pwire FA_out_2488;
  (* register *) pwire FA_out_2489;
  (* register *) pwire FA_out_2490;
  (* register *) pwire FA_out_2491;
  (* register *) pwire FA_out_2492;
  (* register *) pwire FA_out_2493;
  (* register *) pwire FA_out_2494;
  (* register *) pwire FA_out_2495;
  (* register *) pwire FA_out_2496;
  (* register *) pwire FA_out_2497;
  (* register *) pwire FA_out_2498;
  (* register *) pwire FA_out_2499;
  (* register *) pwire FA_out_2500;
  (* register *) pwire FA_out_2501;
  (* register *) pwire FA_out_2502;
  (* register *) pwire FA_out_2503;
  (* register *) pwire FA_out_2504;
  (* register *) pwire FA_out_2505;
  (* register *) pwire FA_out_2506;
  (* register *) pwire FA_out_2507;
  (* register *) pwire FA_out_2508;
  (* register *) pwire FA_out_2509;
  (* register *) pwire FA_out_2510;
  (* register *) pwire FA_out_2511;
  (* register *) pwire FA_out_2512;
  (* register *) pwire FA_out_2513;
  (* register *) pwire FA_out_2514;
  (* register *) pwire FA_out_2515;
  (* register *) pwire FA_out_2516;
  (* register *) pwire FA_out_2517;
  (* register *) pwire FA_out_2518;
  (* register *) pwire FA_out_2519;
  (* register *) pwire FA_out_2520;
  (* register *) pwire FA_out_2521;
  (* register *) pwire FA_out_2522;
  (* register *) pwire FA_out_2523;
  (* register *) pwire FA_out_2524;
  (* register *) pwire FA_out_2525;
  (* register *) pwire FA_out_2526;
  (* register *) pwire FA_out_2527;
  (* register *) pwire FA_out_2528;
  (* register *) pwire FA_out_2529;
  (* register *) pwire FA_out_2530;
  (* register *) pwire FA_out_2531;
  (* register *) pwire FA_out_2532;
  (* register *) pwire FA_out_2533;
  (* register *) pwire FA_out_2534;
  (* register *) pwire FA_out_2535;
  (* register *) pwire FA_out_2536;
  (* register *) pwire FA_out_2537;
  (* register *) pwire FA_out_2538;
  (* register *) pwire FA_out_2539;
  (* register *) pwire FA_out_2540;
  (* register *) pwire FA_out_2541;
  (* register *) pwire FA_out_2542;
  (* register *) pwire FA_out_2543;
  (* register *) pwire FA_out_2544;
  (* register *) pwire FA_out_2545;
  (* register *) pwire FA_out_2546;
  (* register *) pwire FA_out_2547;
  (* register *) pwire FA_out_2548;
  (* register *) pwire FA_out_2549;
  (* register *) pwire FA_out_2550;
  (* register *) pwire FA_out_2551;
  (* register *) pwire FA_out_2552;
  (* register *) pwire FA_out_2553;
  (* register *) pwire FA_out_2554;
  (* register *) pwire FA_out_2555;
  (* register *) pwire FA_out_2556;
  (* register *) pwire FA_out_2557;
  (* register *) pwire FA_out_2558;
  (* register *) pwire FA_out_2559;
  (* register *) pwire FA_out_2560;
  (* register *) pwire FA_out_2561;
  (* register *) pwire FA_out_2562;
  (* register *) pwire FA_out_2563;
  (* register *) pwire FA_out_2564;
  (* register *) pwire FA_out_2565;
  (* register *) pwire FA_out_2566;
  (* register *) pwire FA_out_2567;
  (* register *) pwire FA_out_2568;
  (* register *) pwire FA_out_2569;
  (* register *) pwire FA_out_2570;
  (* register *) pwire FA_out_2571;
  (* register *) pwire FA_out_2572;
  (* register *) pwire FA_out_2573;
  (* register *) pwire FA_out_2574;
  (* register *) pwire FA_out_2575;
  (* register *) pwire FA_out_2576;
  (* register *) pwire FA_out_2577;
  (* register *) pwire FA_out_2578;
  (* register *) pwire FA_out_2579;
  (* register *) pwire FA_out_2580;
  (* register *) pwire FA_out_2581;
  (* register *) pwire FA_out_2582;
  (* register *) pwire FA_out_2583;
  (* register *) pwire FA_out_2584;
  (* register *) pwire FA_out_2585;
  (* register *) pwire FA_out_2586;
  (* register *) pwire FA_out_2587;
  (* register *) pwire FA_out_2588;
  (* register *) pwire FA_out_2589;
  (* register *) pwire FA_out_2590;
  (* register *) pwire FA_out_2591;
  (* register *) pwire FA_out_2592;
  (* register *) pwire FA_out_2593;
  (* register *) pwire FA_out_2594;
  (* register *) pwire FA_out_2595;
  (* register *) pwire FA_out_2596;
  (* register *) pwire FA_out_2597;
  (* register *) pwire FA_out_2598;
  (* register *) pwire FA_out_2599;
  (* register *) pwire FA_out_2600;
  (* register *) pwire FA_out_2601;
  (* register *) pwire FA_out_2602;
  (* register *) pwire FA_out_2603;
  (* register *) pwire FA_out_2604;
  (* register *) pwire FA_out_2605;
  (* register *) pwire FA_out_2606;
  (* register *) pwire FA_out_2607;
  (* register *) pwire FA_out_2608;
  (* register *) pwire FA_out_2609;
  (* register *) pwire FA_out_2610;
  (* register *) pwire FA_out_2611;
  (* register *) pwire FA_out_2612;
  (* register *) pwire FA_out_2613;
  (* register *) pwire FA_out_2614;
  (* register *) pwire FA_out_2615;
  (* register *) pwire FA_out_2616;
  (* register *) pwire FA_out_2617;
  (* register *) pwire FA_out_2618;
  (* register *) pwire FA_out_2619;
  (* register *) pwire FA_out_2620;
  (* register *) pwire FA_out_2621;
  (* register *) pwire FA_out_2622;
  (* register *) pwire FA_out_2623;
  (* register *) pwire FA_out_2624;
  (* register *) pwire FA_out_2625;
  (* register *) pwire FA_out_2626;
  (* register *) pwire FA_out_2627;
  (* register *) pwire FA_out_2628;
  (* register *) pwire FA_out_2629;
  (* register *) pwire FA_out_2630;
  (* register *) pwire FA_out_2631;
  (* register *) pwire FA_out_2632;
  (* register *) pwire FA_out_2633;
  (* register *) pwire FA_out_2634;
  (* register *) pwire FA_out_2635;
  (* register *) pwire FA_out_2636;
  (* register *) pwire FA_out_2637;
  (* register *) pwire FA_out_2638;
  (* register *) pwire FA_out_2639;
  (* register *) pwire FA_out_2640;
  (* register *) pwire FA_out_2641;
  (* register *) pwire FA_out_2642;
  (* register *) pwire FA_out_2643;
  (* register *) pwire FA_out_2644;
  (* register *) pwire FA_out_2645;
  (* register *) pwire FA_out_2646;
  (* register *) pwire FA_out_2647;
  (* register *) pwire FA_out_2648;
  (* register *) pwire FA_out_2649;
  (* register *) pwire FA_out_2650;
  (* register *) pwire FA_out_2651;
  (* register *) pwire FA_out_2652;
  (* register *) pwire FA_out_2653;
  (* register *) pwire FA_out_2654;
  (* register *) pwire FA_out_2655;
  (* register *) pwire FA_out_2656;
  (* register *) pwire FA_out_2657;
  (* register *) pwire FA_out_2658;
  (* register *) pwire FA_out_2659;
  (* register *) pwire FA_out_2660;
  (* register *) pwire FA_out_2661;
  (* register *) pwire FA_out_2662;
  (* register *) pwire FA_out_2663;
  (* register *) pwire FA_out_2664;
  (* register *) pwire FA_out_2665;
  (* register *) pwire FA_out_2666;
  (* register *) pwire FA_out_2667;
  (* register *) pwire FA_out_2668;
  (* register *) pwire FA_out_2669;
  (* register *) pwire FA_out_2670;
  (* register *) pwire FA_out_2671;
  (* register *) pwire FA_out_2672;
  (* register *) pwire FA_out_2673;
  (* register *) pwire FA_out_2674;
  (* register *) pwire FA_out_2675;
  (* register *) pwire FA_out_2676;
  (* register *) pwire FA_out_2677;
  (* register *) pwire FA_out_2678;
  (* register *) pwire FA_out_2679;
  (* register *) pwire FA_out_2680;
  (* register *) pwire FA_out_2681;
  (* register *) pwire FA_out_2682;
  (* register *) pwire FA_out_2683;
  (* register *) pwire FA_out_2684;
  (* register *) pwire FA_out_2685;
  (* register *) pwire FA_out_2686;
  (* register *) pwire FA_out_2687;
  (* register *) pwire FA_out_2688;
  (* register *) pwire FA_out_2689;
  (* register *) pwire FA_out_2690;
  (* register *) pwire FA_out_2691;
  (* register *) pwire FA_out_2692;
  (* register *) pwire FA_out_2693;
  (* register *) pwire FA_out_2694;
  (* register *) pwire FA_out_2695;
  (* register *) pwire FA_out_2696;
  (* register *) pwire FA_out_2697;
  (* register *) pwire FA_out_2698;
  (* register *) pwire FA_out_2699;
  (* register *) pwire FA_out_2700;
  (* register *) pwire FA_out_2701;
  (* register *) pwire FA_out_2702;
  (* register *) pwire FA_out_2703;
  (* register *) pwire FA_out_2704;
  (* register *) pwire FA_out_2705;
  (* register *) pwire FA_out_2706;
  (* register *) pwire FA_out_2707;
  (* register *) pwire FA_out_2708;
  (* register *) pwire FA_out_2709;
  (* register *) pwire FA_out_2710;
  (* register *) pwire FA_out_2711;
  (* register *) pwire FA_out_2712;
  (* register *) pwire FA_out_2713;
  (* register *) pwire FA_out_2714;
  (* register *) pwire FA_out_2715;
  (* register *) pwire FA_out_2716;
  (* register *) pwire FA_out_2717;
  (* register *) pwire FA_out_2718;
  (* register *) pwire FA_out_2719;
  (* register *) pwire FA_out_2720;
  (* register *) pwire FA_out_2721;
  (* register *) pwire FA_out_2722;
  (* register *) pwire FA_out_2723;
  (* register *) pwire FA_out_2724;
  (* register *) pwire FA_out_2725;
  (* register *) pwire FA_out_2726;
  (* register *) pwire FA_out_2727;
  (* register *) pwire FA_out_2728;
  (* register *) pwire FA_out_2729;
  (* register *) pwire FA_out_2730;
  (* register *) pwire FA_out_2731;
  (* register *) pwire FA_out_2732;
  (* register *) pwire FA_out_2733;
  (* register *) pwire FA_out_2734;
  (* register *) pwire FA_out_2735;
  (* register *) pwire FA_out_2736;
  (* register *) pwire FA_out_2737;
  (* register *) pwire FA_out_2738;
  (* register *) pwire FA_out_2739;
  (* register *) pwire FA_out_2740;
  (* register *) pwire FA_out_2741;
  (* register *) pwire FA_out_2742;
  (* register *) pwire FA_out_2743;
  (* register *) pwire FA_out_2744;
  (* register *) pwire FA_out_2745;
  (* register *) pwire FA_out_2746;
  (* register *) pwire FA_out_2747;
  (* register *) pwire FA_out_2748;
  (* register *) pwire FA_out_2749;
  (* register *) pwire FA_out_2750;
  (* register *) pwire FA_out_2751;
  (* register *) pwire FA_out_2752;
  (* register *) pwire FA_out_2753;
  (* register *) pwire FA_out_2754;
  (* register *) pwire FA_out_2755;
  (* register *) pwire FA_out_2756;
  (* register *) pwire FA_out_2757;
  (* register *) pwire FA_out_2758;
  (* register *) pwire FA_out_2759;
  (* register *) pwire FA_out_2760;
  (* register *) pwire FA_out_2761;
  (* register *) pwire FA_out_2762;
  (* register *) pwire FA_out_2763;
  (* register *) pwire FA_out_2764;
  (* register *) pwire FA_out_2765;
  (* register *) pwire FA_out_2766;
  (* register *) pwire FA_out_2767;
  (* register *) pwire FA_out_2768;
  (* register *) pwire FA_out_2769;
  (* register *) pwire FA_out_2770;
  (* register *) pwire FA_out_2771;
  (* register *) pwire FA_out_2772;
  (* register *) pwire FA_out_2773;
  (* register *) pwire FA_out_2774;
  (* register *) pwire FA_out_2775;
  (* register *) pwire FA_out_2776;
  (* register *) pwire FA_out_2777;
  (* register *) pwire FA_out_2778;
  (* register *) pwire FA_out_2779;
  (* register *) pwire FA_out_2780;
  (* register *) pwire FA_out_2781;
  (* register *) pwire FA_out_2782;
  (* register *) pwire FA_out_2783;
  (* register *) pwire FA_out_2784;
  (* register *) pwire FA_out_2785;
  (* register *) pwire FA_out_2786;
  (* register *) pwire FA_out_2787;
  (* register *) pwire FA_out_2788;
  (* register *) pwire FA_out_2789;
  (* register *) pwire FA_out_2790;
  (* register *) pwire FA_out_2791;
  (* register *) pwire FA_out_2792;
  (* register *) pwire FA_out_2793;
  (* register *) pwire FA_out_2794;
  (* register *) pwire FA_out_2795;
  (* register *) pwire FA_out_2796;
  (* register *) pwire FA_out_2797;
  (* register *) pwire FA_out_2798;
  (* register *) pwire FA_out_2799;
  (* register *) pwire FA_out_2800;
  (* register *) pwire FA_out_2801;
  (* register *) pwire FA_out_2802;
  (* register *) pwire FA_out_2803;
  (* register *) pwire FA_out_2804;
  (* register *) pwire FA_out_2805;
  (* register *) pwire FA_out_2806;
  (* register *) pwire FA_out_2807;
  (* register *) pwire FA_out_2808;
  (* register *) pwire FA_out_2809;
  (* register *) pwire FA_out_2810;
  (* register *) pwire FA_out_2811;
  (* register *) pwire FA_out_2812;
  (* register *) pwire FA_out_2813;
  (* register *) pwire FA_out_2814;
  (* register *) pwire FA_out_2815;
  (* register *) pwire FA_out_2816;
  (* register *) pwire FA_out_2817;
  (* register *) pwire FA_out_2818;
  (* register *) pwire FA_out_2819;
  (* register *) pwire FA_out_2820;
  (* register *) pwire FA_out_2821;
  (* register *) pwire FA_out_2822;
  (* register *) pwire FA_out_2823;
  (* register *) pwire FA_out_2824;
  (* register *) pwire FA_out_2825;
  (* register *) pwire FA_out_2826;
  (* register *) pwire FA_out_2827;
  (* register *) pwire FA_out_2828;
  (* register *) pwire FA_out_2829;
  (* register *) pwire FA_out_2830;
  (* register *) pwire FA_out_2831;
  (* register *) pwire FA_out_2832;
  (* register *) pwire FA_out_2833;
  (* register *) pwire FA_out_2834;
  (* register *) pwire FA_out_2835;
  (* register *) pwire FA_out_2836;
  (* register *) pwire FA_out_2837;
  (* register *) pwire FA_out_2838;
  (* register *) pwire FA_out_2839;
  (* register *) pwire FA_out_2840;
  (* register *) pwire FA_out_2841;
  (* register *) pwire FA_out_2842;
  (* register *) pwire FA_out_2843;
  (* register *) pwire FA_out_2844;
  (* register *) pwire FA_out_2845;
  (* register *) pwire FA_out_2846;
  (* register *) pwire FA_out_2847;
  (* register *) pwire FA_out_2848;
  (* register *) pwire FA_out_2849;
  (* register *) pwire FA_out_2850;
  (* register *) pwire FA_out_2851;
  (* register *) pwire FA_out_2852;
  (* register *) pwire FA_out_2853;
  (* register *) pwire FA_out_2854;
  (* register *) pwire FA_out_2855;
  (* register *) pwire FA_out_2856;
  (* register *) pwire FA_out_2857;
  (* register *) pwire FA_out_2858;
  (* register *) pwire FA_out_2859;
  (* register *) pwire FA_out_2860;
  (* register *) pwire FA_out_2861;
  (* register *) pwire FA_out_2862;
  (* register *) pwire FA_out_2863;
  (* register *) pwire FA_out_2864;
  (* register *) pwire FA_out_2865;
  (* register *) pwire FA_out_2866;
  (* register *) pwire FA_out_2867;
  (* register *) pwire FA_out_2868;
  (* register *) pwire FA_out_2869;
  (* register *) pwire FA_out_2870;
  (* register *) pwire FA_out_2871;
  (* register *) pwire FA_out_2872;
  (* register *) pwire FA_out_2873;
  (* register *) pwire FA_out_2874;
  (* register *) pwire FA_out_2875;
  (* register *) pwire FA_out_2876;
  (* register *) pwire FA_out_2877;
  (* register *) pwire FA_out_2878;
  (* register *) pwire FA_out_2879;
  (* register *) pwire FA_out_2880;
  (* register *) pwire FA_out_2881;
  (* register *) pwire FA_out_2882;
  (* register *) pwire FA_out_2883;
  (* register *) pwire FA_out_2884;
  (* register *) pwire FA_out_2885;
  (* register *) pwire FA_out_2886;
  (* register *) pwire FA_out_2887;
  (* register *) pwire FA_out_2888;
  (* register *) pwire FA_out_2889;
  (* register *) pwire FA_out_2890;
  (* register *) pwire FA_out_2891;
  (* register *) pwire FA_out_2892;
  (* register *) pwire FA_out_2893;
  (* register *) pwire FA_out_2894;
  (* register *) pwire FA_out_2895;
  (* register *) pwire FA_out_2896;
  (* register *) pwire FA_out_2897;
  (* register *) pwire FA_out_2898;
  (* register *) pwire FA_out_2899;
  (* register *) pwire FA_out_2900;
  (* register *) pwire FA_out_2901;
  (* register *) pwire FA_out_2902;
  (* register *) pwire FA_out_2903;
  (* register *) pwire FA_out_2904;
  (* register *) pwire FA_out_2905;
  (* register *) pwire FA_out_2906;
  (* register *) pwire FA_out_2907;
  (* register *) pwire FA_out_2908;
  (* register *) pwire FA_out_2909;
  (* register *) pwire FA_out_2910;
  (* register *) pwire FA_out_2911;
  (* register *) pwire FA_out_2912;
  (* register *) pwire FA_out_2913;
  (* register *) pwire FA_out_2914;
  (* register *) pwire FA_out_2915;
  (* register *) pwire FA_out_2916;
  (* register *) pwire FA_out_2917;
  (* register *) pwire FA_out_2918;
  (* register *) pwire FA_out_2919;
  (* register *) pwire FA_out_2920;
  (* register *) pwire FA_out_2921;
  (* register *) pwire FA_out_2922;
  (* register *) pwire FA_out_2923;
  (* register *) pwire FA_out_2924;
  (* register *) pwire FA_out_2925;
  (* register *) pwire FA_out_2926;
  (* register *) pwire FA_out_2927;
  (* register *) pwire FA_out_2928;
  (* register *) pwire FA_out_2929;
  (* register *) pwire FA_out_2930;
  (* register *) pwire FA_out_2931;
  (* register *) pwire FA_out_2932;
  (* register *) pwire FA_out_2933;
  (* register *) pwire FA_out_2934;
  (* register *) pwire FA_out_2935;
  (* register *) pwire FA_out_2936;
  (* register *) pwire FA_out_2937;
  (* register *) pwire FA_out_2938;
  (* register *) pwire FA_out_2939;
  (* register *) pwire FA_out_2940;
  (* register *) pwire FA_out_2941;
  (* register *) pwire FA_out_2942;
  (* register *) pwire FA_out_2943;
  (* register *) pwire FA_out_2944;
  (* register *) pwire FA_out_2945;
  (* register *) pwire FA_out_2946;
  (* register *) pwire FA_out_2947;
  (* register *) pwire FA_out_2948;
  (* register *) pwire FA_out_2949;
  (* register *) pwire FA_out_2950;
  (* register *) pwire FA_out_2951;
  (* register *) pwire FA_out_2952;
  (* register *) pwire FA_out_2953;
  (* register *) pwire FA_out_2954;
  (* register *) pwire FA_out_2955;
  (* register *) pwire FA_out_2956;
  (* register *) pwire FA_out_2957;
  (* register *) pwire FA_out_2958;
  (* register *) pwire FA_out_2959;
  (* register *) pwire FA_out_2960;
  (* register *) pwire FA_out_2961;
  (* register *) pwire FA_out_2962;
  (* register *) pwire FA_out_2963;
  (* register *) pwire FA_out_2964;
  (* register *) pwire FA_out_2965;
  (* register *) pwire FA_out_2966;
  (* register *) pwire FA_out_2967;
  (* register *) pwire FA_out_2968;
  (* register *) pwire FA_out_2969;
  (* register *) pwire FA_out_2970;
  (* register *) pwire FA_out_2971;
  (* register *) pwire FA_out_2972;
  (* register *) pwire FA_out_2973;
  (* register *) pwire FA_out_2974;
  (* register *) pwire FA_out_2975;
  (* register *) pwire FA_out_2976;
  (* register *) pwire FA_out_2977;
  (* register *) pwire FA_out_2978;
  (* register *) pwire FA_out_2979;
  (* register *) pwire FA_out_2980;
  (* register *) pwire FA_out_2981;
  (* register *) pwire FA_out_2982;
  (* register *) pwire FA_out_2983;
  (* register *) pwire FA_out_2984;
  (* register *) pwire FA_out_2985;
  (* register *) pwire FA_out_2986;
  (* register *) pwire FA_out_2987;
  (* register *) pwire FA_out_2988;
  (* register *) pwire FA_out_2989;
  (* register *) pwire FA_out_2990;
  (* register *) pwire FA_out_2991;
  (* register *) pwire FA_out_2992;
  (* register *) pwire FA_out_2993;
  (* register *) pwire FA_out_2994;
  (* register *) pwire FA_out_2995;
  (* register *) pwire FA_out_2996;
  (* register *) pwire FA_out_2997;
  (* register *) pwire FA_out_2998;
  (* register *) pwire FA_out_2999;
  (* register *) pwire FA_out_3000;
  (* register *) pwire FA_out_3001;
  (* register *) pwire FA_out_3002;
  (* register *) pwire FA_out_3003;
  (* register *) pwire FA_out_3004;
  (* register *) pwire FA_out_3005;
  (* register *) pwire FA_out_3006;
  (* register *) pwire FA_out_3007;
  (* register *) pwire FA_out_3008;
  (* register *) pwire FA_out_3009;
  (* register *) pwire FA_out_3010;
  (* register *) pwire FA_out_3011;
  (* register *) pwire FA_out_3012;
  (* register *) pwire FA_out_3013;
  (* register *) pwire FA_out_3014;
  (* register *) pwire FA_out_3015;
  (* register *) pwire FA_out_3016;
  (* register *) pwire FA_out_3017;
  (* register *) pwire FA_out_3018;
  (* register *) pwire FA_out_3019;
  (* register *) pwire FA_out_3020;
  (* register *) pwire FA_out_3021;
  (* register *) pwire FA_out_3022;
  (* register *) pwire FA_out_3023;
  (* register *) pwire FA_out_3024;
  (* register *) pwire FA_out_3025;
  (* register *) pwire FA_out_3026;
  (* register *) pwire FA_out_3027;
  (* register *) pwire FA_out_3028;
  (* register *) pwire FA_out_3029;
  (* register *) pwire FA_out_3030;
  (* register *) pwire FA_out_3031;
  (* register *) pwire FA_out_3032;
  (* register *) pwire FA_out_3033;
  (* register *) pwire FA_out_3034;
  (* register *) pwire FA_out_3035;
  (* register *) pwire FA_out_3036;
  (* register *) pwire FA_out_3037;
  (* register *) pwire FA_out_3038;
  (* register *) pwire FA_out_3039;
  (* register *) pwire FA_out_3040;
  (* register *) pwire FA_out_3041;
  (* register *) pwire FA_out_3042;
  (* register *) pwire FA_out_3043;
  (* register *) pwire FA_out_3044;
  (* register *) pwire FA_out_3045;
  (* register *) pwire FA_out_3046;
  (* register *) pwire FA_out_3047;
  (* register *) pwire FA_out_3048;
  (* register *) pwire FA_out_3049;
  (* register *) pwire FA_out_3050;
  (* register *) pwire FA_out_3051;
  (* register *) pwire FA_out_3052;
  (* register *) pwire FA_out_3053;
  (* register *) pwire FA_out_3054;
  (* register *) pwire FA_out_3055;
  (* register *) pwire FA_out_3056;
  (* register *) pwire FA_out_3057;
  (* register *) pwire FA_out_3058;
  (* register *) pwire FA_out_3059;
  (* register *) pwire FA_out_3060;
  (* register *) pwire FA_out_3061;
  (* register *) pwire FA_out_3062;
  (* register *) pwire FA_out_3063;
  (* register *) pwire FA_out_3064;
  (* register *) pwire FA_out_3065;
  (* register *) pwire FA_out_3066;
  (* register *) pwire FA_out_3067;
  (* register *) pwire FA_out_3068;
  (* register *) pwire FA_out_3069;
  (* register *) pwire FA_out_3070;
  (* register *) pwire FA_out_3071;
  (* register *) pwire FA_out_3072;
  (* register *) pwire FA_out_3073;
  (* register *) pwire FA_out_3074;
  (* register *) pwire FA_out_3075;
  (* register *) pwire FA_out_3076;
  (* register *) pwire FA_out_3077;
  (* register *) pwire FA_out_3078;
  (* register *) pwire FA_out_3079;
  (* register *) pwire FA_out_3080;
  (* register *) pwire FA_out_3081;
  (* register *) pwire FA_out_3082;
  (* register *) pwire FA_out_3083;
  (* register *) pwire FA_out_3084;
  (* register *) pwire FA_out_3085;
  (* register *) pwire FA_out_3086;
  (* register *) pwire FA_out_3087;
  (* register *) pwire FA_out_3088;
  (* register *) pwire FA_out_3089;
  (* register *) pwire FA_out_3090;
  (* register *) pwire FA_out_3091;
  (* register *) pwire FA_out_3092;
  (* register *) pwire FA_out_3093;
  (* register *) pwire FA_out_3094;
  (* register *) pwire FA_out_3095;
  (* register *) pwire FA_out_3096;
  (* register *) pwire FA_out_3097;
  (* register *) pwire FA_out_3098;
  (* register *) pwire FA_out_3099;
  (* register *) pwire FA_out_3100;
  (* register *) pwire FA_out_3101;
  (* register *) pwire FA_out_3102;
  (* register *) pwire FA_out_3103;
  (* register *) pwire FA_out_3104;
  (* register *) pwire FA_out_3105;
  (* register *) pwire FA_out_3106;
  (* register *) pwire FA_out_3107;
  (* register *) pwire FA_out_3108;
  (* register *) pwire FA_out_3109;
  (* register *) pwire FA_out_3110;
  (* register *) pwire FA_out_3111;
  (* register *) pwire FA_out_3112;
  (* register *) pwire FA_out_3113;
  (* register *) pwire FA_out_3114;
  (* register *) pwire FA_out_3115;
  (* register *) pwire FA_out_3116;
  (* register *) pwire FA_out_3117;
  (* register *) pwire FA_out_3118;
  (* register *) pwire FA_out_3119;
  (* register *) pwire FA_out_3120;
  (* register *) pwire FA_out_3121;
  (* register *) pwire FA_out_3122;
  (* register *) pwire FA_out_3123;
  (* register *) pwire FA_out_3124;
  (* register *) pwire FA_out_3125;
  (* register *) pwire FA_out_3126;
  (* register *) pwire FA_out_3127;
  (* register *) pwire FA_out_3128;
  (* register *) pwire FA_out_3129;
  (* register *) pwire FA_out_3130;
  (* register *) pwire FA_out_3131;
  (* register *) pwire FA_out_3132;
  (* register *) pwire FA_out_3133;
  (* register *) pwire FA_out_3134;
  (* register *) pwire FA_out_3135;
  (* register *) pwire FA_out_3136;
  (* register *) pwire FA_out_3137;
  (* register *) pwire FA_out_3138;
  (* register *) pwire FA_out_3139;
  (* register *) pwire FA_out_3140;
  (* register *) pwire FA_out_3141;
  (* register *) pwire FA_out_3142;
  (* register *) pwire FA_out_3143;
  (* register *) pwire FA_out_3144;
  (* register *) pwire FA_out_3145;
  (* register *) pwire FA_out_3146;
  (* register *) pwire FA_out_3147;
  (* register *) pwire FA_out_3148;
  (* register *) pwire FA_out_3149;
  (* register *) pwire FA_out_3150;
  (* register *) pwire FA_out_3151;
  (* register *) pwire FA_out_3152;
  (* register *) pwire FA_out_3153;
  (* register *) pwire FA_out_3154;
  (* register *) pwire FA_out_3155;
  (* register *) pwire FA_out_3156;
  (* register *) pwire FA_out_3157;
  (* register *) pwire FA_out_3158;
  (* register *) pwire FA_out_3159;
  (* register *) pwire FA_out_3160;
  (* register *) pwire FA_out_3161;
  (* register *) pwire FA_out_3162;
  (* register *) pwire FA_out_3163;
  (* register *) pwire FA_out_3164;
  (* register *) pwire FA_out_3165;
  (* register *) pwire FA_out_3166;
  (* register *) pwire FA_out_3167;
  (* register *) pwire FA_out_3168;
  (* register *) pwire FA_out_3169;
  (* register *) pwire FA_out_3170;
  (* register *) pwire FA_out_3171;
  (* register *) pwire FA_out_3172;
  (* register *) pwire FA_out_3173;
  (* register *) pwire FA_out_3174;
  (* register *) pwire FA_out_3175;
  (* register *) pwire FA_out_3176;
  (* register *) pwire FA_out_3177;
  (* register *) pwire FA_out_3178;
  (* register *) pwire FA_out_3179;
  (* register *) pwire FA_out_3180;
  (* register *) pwire FA_out_3181;
  (* register *) pwire FA_out_3182;
  (* register *) pwire FA_out_3183;
  (* register *) pwire FA_out_3184;
  (* register *) pwire FA_out_3185;
  (* register *) pwire FA_out_3186;
  (* register *) pwire FA_out_3187;
  (* register *) pwire FA_out_3188;
  (* register *) pwire FA_out_3189;
  (* register *) pwire FA_out_3190;
  (* register *) pwire FA_out_3191;
  (* register *) pwire FA_out_3192;
  (* register *) pwire FA_out_3193;
  (* register *) pwire FA_out_3194;
  (* register *) pwire FA_out_3195;
  (* register *) pwire FA_out_3196;
  (* register *) pwire FA_out_3197;
  (* register *) pwire FA_out_3198;
  (* register *) pwire FA_out_3199;
  (* register *) pwire FA_out_3200;
  (* register *) pwire FA_out_3201;
  (* register *) pwire FA_out_3202;
  (* register *) pwire FA_out_3203;
  (* register *) pwire FA_out_3204;
  (* register *) pwire FA_out_3205;
  (* register *) pwire FA_out_3206;
  (* register *) pwire FA_out_3207;
  (* register *) pwire FA_out_3208;
  (* register *) pwire FA_out_3209;
  (* register *) pwire FA_out_3210;
  (* register *) pwire FA_out_3211;
  (* register *) pwire FA_out_3212;
  (* register *) pwire FA_out_3213;
  (* register *) pwire FA_out_3214;
  (* register *) pwire FA_out_3215;
  (* register *) pwire FA_out_3216;
  (* register *) pwire FA_out_3217;
  (* register *) pwire FA_out_3218;
  (* register *) pwire FA_out_3219;
  (* register *) pwire FA_out_3220;
  (* register *) pwire FA_out_3221;
  (* register *) pwire FA_out_3222;
  (* register *) pwire FA_out_3223;
  (* register *) pwire FA_out_3224;
  (* register *) pwire FA_out_3225;
  (* register *) pwire FA_out_3226;
  (* register *) pwire FA_out_3227;
  (* register *) pwire FA_out_3228;
  (* register *) pwire FA_out_3229;
  (* register *) pwire FA_out_3230;
  (* register *) pwire FA_out_3231;
  (* register *) pwire FA_out_3232;
  (* register *) pwire FA_out_3233;
  (* register *) pwire FA_out_3234;
  (* register *) pwire FA_out_3235;
  (* register *) pwire FA_out_3236;
  (* register *) pwire FA_out_3237;
  (* register *) pwire FA_out_3238;
  (* register *) pwire FA_out_3239;
  (* register *) pwire FA_out_3240;
  (* register *) pwire FA_out_3241;
  (* register *) pwire FA_out_3242;
  (* register *) pwire FA_out_3243;
  (* register *) pwire FA_out_3244;
  (* register *) pwire FA_out_3245;
  (* register *) pwire FA_out_3246;
  (* register *) pwire FA_out_3247;
  (* register *) pwire FA_out_3248;
  (* register *) pwire FA_out_3249;
  (* register *) pwire FA_out_3250;
  (* register *) pwire FA_out_3251;
  (* register *) pwire FA_out_3252;
  (* register *) pwire FA_out_3253;
  (* register *) pwire FA_out_3254;
  (* register *) pwire FA_out_3255;
  (* register *) pwire FA_out_3256;
  (* register *) pwire FA_out_3257;
  (* register *) pwire FA_out_3258;
  (* register *) pwire FA_out_3259;
  (* register *) pwire FA_out_3260;
  (* register *) pwire FA_out_3261;
  (* register *) pwire FA_out_3262;
  (* register *) pwire FA_out_3263;
  (* register *) pwire FA_out_3264;
  (* register *) pwire FA_out_3265;
  (* register *) pwire FA_out_3266;
  (* register *) pwire FA_out_3267;
  (* register *) pwire FA_out_3268;
  (* register *) pwire FA_out_3269;
  (* register *) pwire FA_out_3270;
  (* register *) pwire FA_out_3271;
  (* register *) pwire FA_out_3272;
  (* register *) pwire FA_out_3273;
  (* register *) pwire FA_out_3274;
  (* register *) pwire FA_out_3275;
  (* register *) pwire FA_out_3276;
  (* register *) pwire FA_out_3277;
  (* register *) pwire FA_out_3278;
  (* register *) pwire FA_out_3279;
  (* register *) pwire FA_out_3280;
  (* register *) pwire FA_out_3281;
  (* register *) pwire FA_out_3282;
  (* register *) pwire FA_out_3283;
  (* register *) pwire FA_out_3284;
  (* register *) pwire FA_out_3285;
  (* register *) pwire FA_out_3286;
  (* register *) pwire FA_out_3287;
  (* register *) pwire FA_out_3288;
  (* register *) pwire FA_out_3289;
  (* register *) pwire FA_out_3290;
  (* register *) pwire FA_out_3291;
  (* register *) pwire FA_out_3292;
  (* register *) pwire FA_out_3293;
  (* register *) pwire FA_out_3294;
  (* register *) pwire FA_out_3295;
  (* register *) pwire FA_out_3296;
  (* register *) pwire FA_out_3297;
  (* register *) pwire FA_out_3298;
  (* register *) pwire FA_out_3299;
  (* register *) pwire FA_out_3300;
  (* register *) pwire FA_out_3301;
  (* register *) pwire FA_out_3302;
  (* register *) pwire FA_out_3303;
  (* register *) pwire FA_out_3304;
  (* register *) pwire FA_out_3305;
  (* register *) pwire FA_out_3306;
  (* register *) pwire FA_out_3307;
  (* register *) pwire FA_out_3308;
  (* register *) pwire FA_out_3309;
  (* register *) pwire FA_out_3310;
  (* register *) pwire FA_out_3311;
  (* register *) pwire FA_out_3312;
  (* register *) pwire FA_out_3313;
  (* register *) pwire FA_out_3314;
  (* register *) pwire FA_out_3315;
  (* register *) pwire FA_out_3316;
  (* register *) pwire FA_out_3317;
  (* register *) pwire FA_out_3318;
  (* register *) pwire FA_out_3319;
  (* register *) pwire FA_out_3320;
  (* register *) pwire FA_out_3321;
  (* register *) pwire FA_out_3322;
  (* register *) pwire FA_out_3323;
  (* register *) pwire FA_out_3324;
  (* register *) pwire FA_out_3325;
  (* register *) pwire FA_out_3326;
  (* register *) pwire FA_out_3327;
  (* register *) pwire FA_out_3328;
  (* register *) pwire FA_out_3329;
  (* register *) pwire FA_out_3330;
  (* register *) pwire FA_out_3331;
  (* register *) pwire FA_out_3332;
  (* register *) pwire FA_out_3333;
  (* register *) pwire FA_out_3334;
  (* register *) pwire FA_out_3335;
  (* register *) pwire FA_out_3336;
  (* register *) pwire FA_out_3337;
  (* register *) pwire FA_out_3338;
  (* register *) pwire FA_out_3339;
  (* register *) pwire FA_out_3340;
  (* register *) pwire FA_out_3341;
  (* register *) pwire FA_out_3342;
  (* register *) pwire FA_out_3343;
  (* register *) pwire FA_out_3344;
  (* register *) pwire FA_out_3345;
  (* register *) pwire FA_out_3346;
  (* register *) pwire FA_out_3347;
  (* register *) pwire FA_out_3348;
  (* register *) pwire FA_out_3349;
  (* register *) pwire FA_out_3350;
  (* register *) pwire FA_out_3351;
  (* register *) pwire FA_out_3352;
  (* register *) pwire FA_out_3353;
  (* register *) pwire FA_out_3354;
  (* register *) pwire FA_out_3355;
  (* register *) pwire FA_out_3356;
  (* register *) pwire FA_out_3357;
  (* register *) pwire FA_out_3358;
  (* register *) pwire FA_out_3359;
  (* register *) pwire FA_out_3360;
  (* register *) pwire FA_out_3361;
  (* register *) pwire FA_out_3362;
  (* register *) pwire FA_out_3363;
  (* register *) pwire FA_out_3364;
  (* register *) pwire FA_out_3365;
  (* register *) pwire FA_out_3366;
  (* register *) pwire FA_out_3367;
  (* register *) pwire FA_out_3368;
  (* register *) pwire FA_out_3369;
  (* register *) pwire FA_out_3370;
  (* register *) pwire FA_out_3371;
  (* register *) pwire FA_out_3372;
  (* register *) pwire FA_out_3373;
  (* register *) pwire FA_out_3374;
  (* register *) pwire FA_out_3375;
  (* register *) pwire FA_out_3376;
  (* register *) pwire FA_out_3377;
  (* register *) pwire FA_out_3378;
  (* register *) pwire FA_out_3379;
  (* register *) pwire FA_out_3380;
  (* register *) pwire FA_out_3381;
  (* register *) pwire FA_out_3382;
  (* register *) pwire FA_out_3383;
  (* register *) pwire FA_out_3384;
  (* register *) pwire FA_out_3385;
  (* register *) pwire FA_out_3386;
  (* register *) pwire FA_out_3387;
  (* register *) pwire FA_out_3388;
  (* register *) pwire FA_out_3389;
  (* register *) pwire FA_out_3390;
  (* register *) pwire FA_out_3391;
  (* register *) pwire FA_out_3392;
  (* register *) pwire FA_out_3393;
  (* register *) pwire FA_out_3394;
  (* register *) pwire FA_out_3395;
  (* register *) pwire FA_out_3396;
  (* register *) pwire FA_out_3397;
  (* register *) pwire FA_out_3398;
  (* register *) pwire FA_out_3399;
  (* register *) pwire FA_out_3400;
  (* register *) pwire FA_out_3401;
  (* register *) pwire FA_out_3402;
  (* register *) pwire FA_out_3403;
  (* register *) pwire FA_out_3404;
  (* register *) pwire FA_out_3405;
  (* register *) pwire FA_out_3406;
  (* register *) pwire FA_out_3407;
  (* register *) pwire FA_out_3408;
  (* register *) pwire FA_out_3409;
  (* register *) pwire FA_out_3410;
  (* register *) pwire FA_out_3411;
  (* register *) pwire FA_out_3412;
  (* register *) pwire FA_out_3413;
  (* register *) pwire FA_out_3414;
  (* register *) pwire FA_out_3415;
  (* register *) pwire FA_out_3416;
  (* register *) pwire FA_out_3417;
  (* register *) pwire FA_out_3418;
  (* register *) pwire FA_out_3419;
  (* register *) pwire FA_out_3420;
  (* register *) pwire FA_out_3421;
  (* register *) pwire FA_out_3422;
  (* register *) pwire FA_out_3423;
  (* register *) pwire FA_out_3424;
  (* register *) pwire FA_out_3425;
  (* register *) pwire FA_out_3426;
  (* register *) pwire FA_out_3427;
  (* register *) pwire FA_out_3428;
  (* register *) pwire FA_out_3429;
  (* register *) pwire FA_out_3430;
  (* register *) pwire FA_out_3431;
  (* register *) pwire FA_out_3432;
  (* register *) pwire FA_out_3433;
  (* register *) pwire FA_out_3434;
  (* register *) pwire FA_out_3435;
  (* register *) pwire FA_out_3436;
  (* register *) pwire FA_out_3437;
  (* register *) pwire FA_out_3438;
  (* register *) pwire FA_out_3439;
  (* register *) pwire FA_out_3440;
  (* register *) pwire FA_out_3441;
  (* register *) pwire FA_out_3442;
  (* register *) pwire FA_out_3443;
  (* register *) pwire FA_out_3444;
  (* register *) pwire FA_out_3445;
  (* register *) pwire FA_out_3446;
  (* register *) pwire FA_out_3447;
  (* register *) pwire FA_out_3448;
  (* register *) pwire FA_out_3449;
  (* register *) pwire FA_out_3450;
  (* register *) pwire FA_out_3451;
  (* register *) pwire FA_out_3452;
  (* register *) pwire FA_out_3453;
  (* register *) pwire FA_out_3454;
  (* register *) pwire FA_out_3455;
  (* register *) pwire FA_out_3456;
  (* register *) pwire FA_out_3457;
  (* register *) pwire FA_out_3458;
  (* register *) pwire FA_out_3459;
  (* register *) pwire FA_out_3460;
  (* register *) pwire FA_out_3461;
  (* register *) pwire FA_out_3462;
  (* register *) pwire FA_out_3463;
  (* register *) pwire FA_out_3464;
  (* register *) pwire FA_out_3465;
  (* register *) pwire FA_out_3466;
  (* register *) pwire FA_out_3467;
  (* register *) pwire FA_out_3468;
  (* register *) pwire FA_out_3469;
  (* register *) pwire FA_out_3470;
  (* register *) pwire FA_out_3471;
  (* register *) pwire FA_out_3472;
  (* register *) pwire FA_out_3473;
  (* register *) pwire FA_out_3474;
  (* register *) pwire FA_out_3475;
  (* register *) pwire FA_out_3476;
  (* register *) pwire FA_out_3477;
  (* register *) pwire FA_out_3478;
  (* register *) pwire FA_out_3479;
  (* register *) pwire FA_out_3480;
  (* register *) pwire FA_out_3481;
  (* register *) pwire FA_out_3482;
  (* register *) pwire FA_out_3483;
  (* register *) pwire FA_out_3484;
  (* register *) pwire FA_out_3485;
  (* register *) pwire FA_out_3486;
  (* register *) pwire FA_out_3487;
  (* register *) pwire FA_out_3488;
  (* register *) pwire FA_out_3489;
  (* register *) pwire FA_out_3490;
  (* register *) pwire FA_out_3491;
  (* register *) pwire FA_out_3492;
  (* register *) pwire FA_out_3493;
  (* register *) pwire FA_out_3494;
  (* register *) pwire FA_out_3495;
  (* register *) pwire FA_out_3496;
  (* register *) pwire FA_out_3497;
  (* register *) pwire FA_out_3498;
  (* register *) pwire FA_out_3499;
  (* register *) pwire FA_out_3500;
  (* register *) pwire FA_out_3501;
  (* register *) pwire FA_out_3502;
  (* register *) pwire FA_out_3503;
  (* register *) pwire FA_out_3504;
  (* register *) pwire FA_out_3505;
  (* register *) pwire FA_out_3506;
  (* register *) pwire FA_out_3507;
  (* register *) pwire FA_out_3508;
  (* register *) pwire FA_out_3509;
  (* register *) pwire FA_out_3510;
  (* register *) pwire FA_out_3511;
  (* register *) pwire FA_out_3512;
  (* register *) pwire FA_out_3513;
  (* register *) pwire FA_out_3514;
  (* register *) pwire FA_out_3515;
  (* register *) pwire FA_out_3516;
  (* register *) pwire FA_out_3517;
  (* register *) pwire FA_out_3518;
  (* register *) pwire FA_out_3519;
  (* register *) pwire FA_out_3520;
  (* register *) pwire FA_out_3521;
  (* register *) pwire FA_out_3522;
  (* register *) pwire FA_out_3523;
  (* register *) pwire FA_out_3524;
  (* register *) pwire FA_out_3525;
  (* register *) pwire FA_out_3526;
  (* register *) pwire FA_out_3527;
  (* register *) pwire FA_out_3528;
  (* register *) pwire FA_out_3529;
  (* register *) pwire FA_out_3530;
  (* register *) pwire FA_out_3531;
  (* register *) pwire FA_out_3532;
  (* register *) pwire FA_out_3533;
  (* register *) pwire FA_out_3534;
  (* register *) pwire FA_out_3535;
  (* register *) pwire FA_out_3536;
  (* register *) pwire FA_out_3537;
  (* register *) pwire FA_out_3538;
  (* register *) pwire FA_out_3539;
  (* register *) pwire FA_out_3540;
  (* register *) pwire FA_out_3541;
  (* register *) pwire FA_out_3542;
  (* register *) pwire FA_out_3543;
  (* register *) pwire FA_out_3544;
  (* register *) pwire FA_out_3545;
  (* register *) pwire FA_out_3546;
  (* register *) pwire FA_out_3547;
  (* register *) pwire FA_out_3548;
  (* register *) pwire FA_out_3549;
  (* register *) pwire FA_out_3550;
  (* register *) pwire FA_out_3551;
  (* register *) pwire FA_out_3552;
  (* register *) pwire FA_out_3553;
  (* register *) pwire FA_out_3554;
  (* register *) pwire FA_out_3555;
  (* register *) pwire FA_out_3556;
  (* register *) pwire FA_out_3557;
  (* register *) pwire FA_out_3558;
  (* register *) pwire FA_out_3559;
  (* register *) pwire FA_out_3560;
  (* register *) pwire FA_out_3561;
  (* register *) pwire FA_out_3562;
  (* register *) pwire FA_out_3563;
  (* register *) pwire FA_out_3564;
  (* register *) pwire FA_out_3565;
  (* register *) pwire FA_out_3566;
  (* register *) pwire FA_out_3567;
  (* register *) pwire FA_out_3568;
  (* register *) pwire FA_out_3569;
  (* register *) pwire FA_out_3570;
  (* register *) pwire FA_out_3571;
  (* register *) pwire FA_out_3572;
  (* register *) pwire FA_out_3573;
  (* register *) pwire FA_out_3574;
  (* register *) pwire FA_out_3575;
  (* register *) pwire FA_out_3576;
  (* register *) pwire FA_out_3577;
  (* register *) pwire FA_out_3578;
  (* register *) pwire FA_out_3579;
  (* register *) pwire FA_out_3580;
  (* register *) pwire FA_out_3581;
  (* register *) pwire FA_out_3582;
  (* register *) pwire FA_out_3583;
  (* register *) pwire FA_out_3584;
  (* register *) pwire FA_out_3585;
  (* register *) pwire FA_out_3586;
  (* register *) pwire FA_out_3587;
  (* register *) pwire FA_out_3588;
  (* register *) pwire FA_out_3589;
  (* register *) pwire FA_out_3590;
  (* register *) pwire FA_out_3591;
  (* register *) pwire FA_out_3592;
  (* register *) pwire FA_out_3593;
  (* register *) pwire FA_out_3594;
  (* register *) pwire FA_out_3595;
  (* register *) pwire FA_out_3596;
  (* register *) pwire FA_out_3597;
  (* register *) pwire FA_out_3598;
  (* register *) pwire FA_out_3599;
  (* register *) pwire FA_out_3600;
  (* register *) pwire FA_out_3601;
  (* register *) pwire FA_out_3602;
  (* register *) pwire FA_out_3603;
  (* register *) pwire FA_out_3604;
  (* register *) pwire FA_out_3605;
  (* register *) pwire FA_out_3606;
  (* register *) pwire FA_out_3607;
  (* register *) pwire FA_out_3608;
  (* register *) pwire FA_out_3609;
  (* register *) pwire FA_out_3610;
  (* register *) pwire FA_out_3611;
  (* register *) pwire FA_out_3612;
  (* register *) pwire FA_out_3613;
  (* register *) pwire FA_out_3614;
  (* register *) pwire FA_out_3615;
  (* register *) pwire FA_out_3616;
  (* register *) pwire FA_out_3617;
  (* register *) pwire FA_out_3618;
  (* register *) pwire FA_out_3619;
  (* register *) pwire FA_out_3620;
  (* register *) pwire FA_out_3621;
  (* register *) pwire FA_out_3622;
  (* register *) pwire FA_out_3623;
  (* register *) pwire FA_out_3624;
  (* register *) pwire FA_out_3625;
  (* register *) pwire FA_out_3626;
  (* register *) pwire FA_out_3627;
  (* register *) pwire FA_out_3628;
  (* register *) pwire FA_out_3629;
  (* register *) pwire FA_out_3630;
  (* register *) pwire FA_out_3631;
  (* register *) pwire FA_out_3632;
  (* register *) pwire FA_out_3633;
  (* register *) pwire FA_out_3634;
  (* register *) pwire FA_out_3635;
  (* register *) pwire FA_out_3636;
  (* register *) pwire FA_out_3637;
  (* register *) pwire FA_out_3638;
  (* register *) pwire FA_out_3639;
  (* register *) pwire FA_out_3640;
  (* register *) pwire FA_out_3641;
  (* register *) pwire FA_out_3642;
  (* register *) pwire FA_out_3643;
  (* register *) pwire FA_out_3644;
  (* register *) pwire FA_out_3645;
  (* register *) pwire FA_out_3646;
  (* register *) pwire FA_out_3647;
  (* register *) pwire FA_out_3648;
  (* register *) pwire FA_out_3649;
  (* register *) pwire FA_out_3650;
  (* register *) pwire FA_out_3651;
  (* register *) pwire FA_out_3652;
  (* register *) pwire FA_out_3653;
  (* register *) pwire FA_out_3654;
  (* register *) pwire FA_out_3655;
  (* register *) pwire FA_out_3656;
  (* register *) pwire FA_out_3657;
  (* register *) pwire FA_out_3658;
  (* register *) pwire FA_out_3659;
  (* register *) pwire FA_out_3660;
  (* register *) pwire FA_out_3661;
  (* register *) pwire FA_out_3662;
  (* register *) pwire FA_out_3663;
  (* register *) pwire FA_out_3664;
  (* register *) pwire FA_out_3665;
  (* register *) pwire FA_out_3666;
  (* register *) pwire FA_out_3667;
  (* register *) pwire FA_out_3668;
  (* register *) pwire FA_out_3669;
  (* register *) pwire FA_out_3670;
  (* register *) pwire FA_out_3671;
  (* register *) pwire FA_out_3672;
  (* register *) pwire FA_out_3673;
  (* register *) pwire FA_out_3674;
  (* register *) pwire FA_out_3675;
  (* register *) pwire FA_out_3676;
  (* register *) pwire FA_out_3677;
  (* register *) pwire FA_out_3678;
  (* register *) pwire FA_out_3679;
  (* register *) pwire FA_out_3680;
  (* register *) pwire FA_out_3681;
  (* register *) pwire FA_out_3682;
  (* register *) pwire FA_out_3683;
  (* register *) pwire FA_out_3684;
  (* register *) pwire FA_out_3685;
  (* register *) pwire FA_out_3686;
  (* register *) pwire FA_out_3687;
  (* register *) pwire FA_out_3688;
  (* register *) pwire FA_out_3689;
  (* register *) pwire FA_out_3690;
  (* register *) pwire FA_out_3691;
  (* register *) pwire FA_out_3692;
  (* register *) pwire FA_out_3693;
  (* register *) pwire FA_out_3694;
  (* register *) pwire FA_out_3695;
  (* register *) pwire FA_out_3696;
  (* register *) pwire FA_out_3697;
  (* register *) pwire FA_out_3698;
  (* register *) pwire FA_out_3699;
  (* register *) pwire FA_out_3700;
  (* register *) pwire FA_out_3701;
  (* register *) pwire FA_out_3702;
  (* register *) pwire FA_out_3703;
  (* register *) pwire FA_out_3704;
  (* register *) pwire FA_out_3705;
  (* register *) pwire FA_out_3706;
  (* register *) pwire FA_out_3707;
  (* register *) pwire FA_out_3708;
  (* register *) pwire FA_out_3709;
  (* register *) pwire FA_out_3710;
  (* register *) pwire FA_out_3711;
  (* register *) pwire FA_out_3712;
  (* register *) pwire FA_out_3713;
  (* register *) pwire FA_out_3714;
  (* register *) pwire FA_out_3715;
  (* register *) pwire FA_out_3716;
  (* register *) pwire FA_out_3717;
  (* register *) pwire FA_out_3718;
  (* register *) pwire FA_out_3719;
  (* register *) pwire FA_out_3720;
  (* register *) pwire FA_out_3721;
  (* register *) pwire FA_out_3722;
  (* register *) pwire FA_out_3723;
  (* register *) pwire FA_out_3724;
  (* register *) pwire FA_out_3725;
  (* register *) pwire FA_out_3726;
  (* register *) pwire FA_out_3727;
  (* register *) pwire FA_out_3728;
  (* register *) pwire FA_out_3729;
  (* register *) pwire FA_out_3730;
  (* register *) pwire FA_out_3731;
  (* register *) pwire FA_out_3732;
  (* register *) pwire FA_out_3733;
  (* register *) pwire FA_out_3734;
  (* register *) pwire FA_out_3735;
  (* register *) pwire FA_out_3736;
  (* register *) pwire FA_out_3737;
  (* register *) pwire FA_out_3738;
  (* register *) pwire FA_out_3739;
  (* register *) pwire FA_out_3740;
  (* register *) pwire FA_out_3741;
  (* register *) pwire FA_out_3742;
  (* register *) pwire FA_out_3743;
  (* register *) pwire FA_out_3744;
  (* register *) pwire FA_out_3745;
  (* register *) pwire FA_out_3746;
  (* register *) pwire FA_out_3747;
  (* register *) pwire FA_out_3748;
  (* register *) pwire FA_out_3749;
  (* register *) pwire FA_out_3750;
  (* register *) pwire FA_out_3751;
  (* register *) pwire FA_out_3752;
  (* register *) pwire FA_out_3753;
  (* register *) pwire FA_out_3754;
  (* register *) pwire FA_out_3755;
  (* register *) pwire FA_out_3756;
  (* register *) pwire FA_out_3757;
  (* register *) pwire FA_out_3758;
  (* register *) pwire FA_out_3759;
  (* register *) pwire FA_out_3760;
  (* register *) pwire FA_out_3761;
  (* register *) pwire FA_out_3762;
  (* register *) pwire FA_out_3763;
  (* register *) pwire FA_out_3764;
  (* register *) pwire FA_out_3765;
  (* register *) pwire FA_out_3766;
  (* register *) pwire FA_out_3767;
  (* register *) pwire FA_out_3768;
  (* register *) pwire FA_out_3769;
  (* register *) pwire FA_out_3770;
  (* register *) pwire FA_out_3771;
  (* register *) pwire FA_out_3772;
  (* register *) pwire FA_out_3773;
  (* register *) pwire FA_out_3774;
  (* register *) pwire FA_out_3775;
  (* register *) pwire FA_out_3776;
  (* register *) pwire FA_out_3777;
  (* register *) pwire FA_out_3778;
  (* register *) pwire FA_out_3779;
  (* register *) pwire FA_out_3780;
  (* register *) pwire FA_out_3781;
  (* register *) pwire FA_out_3782;
  (* register *) pwire FA_out_3783;
  (* register *) pwire FA_out_3784;
  (* register *) pwire FA_out_3785;
  (* register *) pwire FA_out_3786;
  (* register *) pwire FA_out_3787;
  (* register *) pwire FA_out_3788;
  (* register *) pwire FA_out_3789;
  (* register *) pwire FA_out_3790;
  (* register *) pwire FA_out_3791;
  (* register *) pwire FA_out_3792;
  (* register *) pwire FA_out_3793;
  (* register *) pwire FA_out_3794;
  (* register *) pwire FA_out_3795;
  (* register *) pwire FA_out_3796;
  (* register *) pwire FA_out_3797;
  (* register *) pwire FA_out_3798;
  (* register *) pwire FA_out_3799;
  (* register *) pwire FA_out_3800;
  (* register *) pwire FA_out_3801;
  (* register *) pwire FA_out_3802;
  (* register *) pwire FA_out_3803;
  (* register *) pwire FA_out_3804;
  (* register *) pwire FA_out_3805;
  (* register *) pwire FA_out_3806;
  (* register *) pwire FA_out_3807;
  (* register *) pwire FA_out_3808;
  (* register *) pwire FA_out_3809;
  (* register *) pwire FA_out_3810;
  (* register *) pwire FA_out_3811;
  (* register *) pwire FA_out_3812;
  (* register *) pwire FA_out_3813;
  (* register *) pwire FA_out_3814;
  (* register *) pwire FA_out_3815;
  (* register *) pwire FA_out_3816;
  (* register *) pwire FA_out_3817;
  (* register *) pwire FA_out_3818;
  (* register *) pwire FA_out_3819;
  (* register *) pwire FA_out_3820;
  (* register *) pwire FA_out_3821;
  (* register *) pwire FA_out_3822;
  (* register *) pwire FA_out_3823;
  (* register *) pwire FA_out_3824;
  (* register *) pwire FA_out_3825;
  (* register *) pwire FA_out_3826;
  (* register *) pwire FA_out_3827;
  (* register *) pwire FA_out_3828;
  (* register *) pwire FA_out_3829;
  (* register *) pwire FA_out_3830;
  (* register *) pwire FA_out_3831;
  (* register *) pwire FA_out_3832;
  (* register *) pwire FA_out_3833;
  (* register *) pwire FA_out_3834;
  (* register *) pwire FA_out_3835;
  (* register *) pwire FA_out_3836;
  (* register *) pwire FA_out_3837;
  (* register *) pwire FA_out_3838;
  (* register *) pwire FA_out_3839;
  (* register *) pwire FA_out_3840;
  (* register *) pwire FA_out_3841;
  (* register *) pwire FA_out_3842;
  (* register *) pwire FA_out_3843;
  (* register *) pwire FA_out_3844;
  (* register *) pwire FA_out_3845;
  (* register *) pwire FA_cout_0;
  (* register *) pwire FA_cout_1;
  (* register *) pwire FA_cout_2;
  (* register *) pwire FA_cout_3;
  (* register *) pwire FA_cout_4;
  (* register *) pwire FA_cout_5;
  (* register *) pwire FA_cout_6;
  (* register *) pwire FA_cout_7;
  (* register *) pwire FA_cout_8;
  (* register *) pwire FA_cout_9;
  (* register *) pwire FA_cout_10;
  (* register *) pwire FA_cout_11;
  (* register *) pwire FA_cout_12;
  (* register *) pwire FA_cout_13;
  (* register *) pwire FA_cout_14;
  (* register *) pwire FA_cout_15;
  (* register *) pwire FA_cout_16;
  (* register *) pwire FA_cout_17;
  (* register *) pwire FA_cout_18;
  (* register *) pwire FA_cout_19;
  (* register *) pwire FA_cout_20;
  (* register *) pwire FA_cout_21;
  (* register *) pwire FA_cout_22;
  (* register *) pwire FA_cout_23;
  (* register *) pwire FA_cout_24;
  (* register *) pwire FA_cout_25;
  (* register *) pwire FA_cout_26;
  (* register *) pwire FA_cout_27;
  (* register *) pwire FA_cout_28;
  (* register *) pwire FA_cout_29;
  (* register *) pwire FA_cout_30;
  (* register *) pwire FA_cout_31;
  (* register *) pwire FA_cout_32;
  (* register *) pwire FA_cout_33;
  (* register *) pwire FA_cout_34;
  (* register *) pwire FA_cout_35;
  (* register *) pwire FA_cout_36;
  (* register *) pwire FA_cout_37;
  (* register *) pwire FA_cout_38;
  (* register *) pwire FA_cout_39;
  (* register *) pwire FA_cout_40;
  (* register *) pwire FA_cout_41;
  (* register *) pwire FA_cout_42;
  (* register *) pwire FA_cout_43;
  (* register *) pwire FA_cout_44;
  (* register *) pwire FA_cout_45;
  (* register *) pwire FA_cout_46;
  (* register *) pwire FA_cout_47;
  (* register *) pwire FA_cout_48;
  (* register *) pwire FA_cout_49;
  (* register *) pwire FA_cout_50;
  (* register *) pwire FA_cout_51;
  (* register *) pwire FA_cout_52;
  (* register *) pwire FA_cout_53;
  (* register *) pwire FA_cout_54;
  (* register *) pwire FA_cout_55;
  (* register *) pwire FA_cout_56;
  (* register *) pwire FA_cout_57;
  (* register *) pwire FA_cout_58;
  (* register *) pwire FA_cout_59;
  (* register *) pwire FA_cout_60;
  (* register *) pwire FA_cout_61;
  (* register *) pwire FA_cout_62;
  (* register *) pwire FA_cout_63;
  (* register *) pwire FA_cout_64;
  (* register *) pwire FA_cout_65;
  (* register *) pwire FA_cout_66;
  (* register *) pwire FA_cout_67;
  (* register *) pwire FA_cout_68;
  (* register *) pwire FA_cout_69;
  (* register *) pwire FA_cout_70;
  (* register *) pwire FA_cout_71;
  (* register *) pwire FA_cout_72;
  (* register *) pwire FA_cout_73;
  (* register *) pwire FA_cout_74;
  (* register *) pwire FA_cout_75;
  (* register *) pwire FA_cout_76;
  (* register *) pwire FA_cout_77;
  (* register *) pwire FA_cout_78;
  (* register *) pwire FA_cout_79;
  (* register *) pwire FA_cout_80;
  (* register *) pwire FA_cout_81;
  (* register *) pwire FA_cout_82;
  (* register *) pwire FA_cout_83;
  (* register *) pwire FA_cout_84;
  (* register *) pwire FA_cout_85;
  (* register *) pwire FA_cout_86;
  (* register *) pwire FA_cout_87;
  (* register *) pwire FA_cout_88;
  (* register *) pwire FA_cout_89;
  (* register *) pwire FA_cout_90;
  (* register *) pwire FA_cout_91;
  (* register *) pwire FA_cout_92;
  (* register *) pwire FA_cout_93;
  (* register *) pwire FA_cout_94;
  (* register *) pwire FA_cout_95;
  (* register *) pwire FA_cout_96;
  (* register *) pwire FA_cout_97;
  (* register *) pwire FA_cout_98;
  (* register *) pwire FA_cout_99;
  (* register *) pwire FA_cout_100;
  (* register *) pwire FA_cout_101;
  (* register *) pwire FA_cout_102;
  (* register *) pwire FA_cout_103;
  (* register *) pwire FA_cout_104;
  (* register *) pwire FA_cout_105;
  (* register *) pwire FA_cout_106;
  (* register *) pwire FA_cout_107;
  (* register *) pwire FA_cout_108;
  (* register *) pwire FA_cout_109;
  (* register *) pwire FA_cout_110;
  (* register *) pwire FA_cout_111;
  (* register *) pwire FA_cout_112;
  (* register *) pwire FA_cout_113;
  (* register *) pwire FA_cout_114;
  (* register *) pwire FA_cout_115;
  (* register *) pwire FA_cout_116;
  (* register *) pwire FA_cout_117;
  (* register *) pwire FA_cout_118;
  (* register *) pwire FA_cout_119;
  (* register *) pwire FA_cout_120;
  (* register *) pwire FA_cout_121;
  (* register *) pwire FA_cout_122;
  (* register *) pwire FA_cout_123;
  (* register *) pwire FA_cout_124;
  (* register *) pwire FA_cout_125;
  (* register *) pwire FA_cout_126;
  (* register *) pwire FA_cout_127;
  (* register *) pwire FA_cout_128;
  (* register *) pwire FA_cout_129;
  (* register *) pwire FA_cout_130;
  (* register *) pwire FA_cout_131;
  (* register *) pwire FA_cout_132;
  (* register *) pwire FA_cout_133;
  (* register *) pwire FA_cout_134;
  (* register *) pwire FA_cout_135;
  (* register *) pwire FA_cout_136;
  (* register *) pwire FA_cout_137;
  (* register *) pwire FA_cout_138;
  (* register *) pwire FA_cout_139;
  (* register *) pwire FA_cout_140;
  (* register *) pwire FA_cout_141;
  (* register *) pwire FA_cout_142;
  (* register *) pwire FA_cout_143;
  (* register *) pwire FA_cout_144;
  (* register *) pwire FA_cout_145;
  (* register *) pwire FA_cout_146;
  (* register *) pwire FA_cout_147;
  (* register *) pwire FA_cout_148;
  (* register *) pwire FA_cout_149;
  (* register *) pwire FA_cout_150;
  (* register *) pwire FA_cout_151;
  (* register *) pwire FA_cout_152;
  (* register *) pwire FA_cout_153;
  (* register *) pwire FA_cout_154;
  (* register *) pwire FA_cout_155;
  (* register *) pwire FA_cout_156;
  (* register *) pwire FA_cout_157;
  (* register *) pwire FA_cout_158;
  (* register *) pwire FA_cout_159;
  (* register *) pwire FA_cout_160;
  (* register *) pwire FA_cout_161;
  (* register *) pwire FA_cout_162;
  (* register *) pwire FA_cout_163;
  (* register *) pwire FA_cout_164;
  (* register *) pwire FA_cout_165;
  (* register *) pwire FA_cout_166;
  (* register *) pwire FA_cout_167;
  (* register *) pwire FA_cout_168;
  (* register *) pwire FA_cout_169;
  (* register *) pwire FA_cout_170;
  (* register *) pwire FA_cout_171;
  (* register *) pwire FA_cout_172;
  (* register *) pwire FA_cout_173;
  (* register *) pwire FA_cout_174;
  (* register *) pwire FA_cout_175;
  (* register *) pwire FA_cout_176;
  (* register *) pwire FA_cout_177;
  (* register *) pwire FA_cout_178;
  (* register *) pwire FA_cout_179;
  (* register *) pwire FA_cout_180;
  (* register *) pwire FA_cout_181;
  (* register *) pwire FA_cout_182;
  (* register *) pwire FA_cout_183;
  (* register *) pwire FA_cout_184;
  (* register *) pwire FA_cout_185;
  (* register *) pwire FA_cout_186;
  (* register *) pwire FA_cout_187;
  (* register *) pwire FA_cout_188;
  (* register *) pwire FA_cout_189;
  (* register *) pwire FA_cout_190;
  (* register *) pwire FA_cout_191;
  (* register *) pwire FA_cout_192;
  (* register *) pwire FA_cout_193;
  (* register *) pwire FA_cout_194;
  (* register *) pwire FA_cout_195;
  (* register *) pwire FA_cout_196;
  (* register *) pwire FA_cout_197;
  (* register *) pwire FA_cout_198;
  (* register *) pwire FA_cout_199;
  (* register *) pwire FA_cout_200;
  (* register *) pwire FA_cout_201;
  (* register *) pwire FA_cout_202;
  (* register *) pwire FA_cout_203;
  (* register *) pwire FA_cout_204;
  (* register *) pwire FA_cout_205;
  (* register *) pwire FA_cout_206;
  (* register *) pwire FA_cout_207;
  (* register *) pwire FA_cout_208;
  (* register *) pwire FA_cout_209;
  (* register *) pwire FA_cout_210;
  (* register *) pwire FA_cout_211;
  (* register *) pwire FA_cout_212;
  (* register *) pwire FA_cout_213;
  (* register *) pwire FA_cout_214;
  (* register *) pwire FA_cout_215;
  (* register *) pwire FA_cout_216;
  (* register *) pwire FA_cout_217;
  (* register *) pwire FA_cout_218;
  (* register *) pwire FA_cout_219;
  (* register *) pwire FA_cout_220;
  (* register *) pwire FA_cout_221;
  (* register *) pwire FA_cout_222;
  (* register *) pwire FA_cout_223;
  (* register *) pwire FA_cout_224;
  (* register *) pwire FA_cout_225;
  (* register *) pwire FA_cout_226;
  (* register *) pwire FA_cout_227;
  (* register *) pwire FA_cout_228;
  (* register *) pwire FA_cout_229;
  (* register *) pwire FA_cout_230;
  (* register *) pwire FA_cout_231;
  (* register *) pwire FA_cout_232;
  (* register *) pwire FA_cout_233;
  (* register *) pwire FA_cout_234;
  (* register *) pwire FA_cout_235;
  (* register *) pwire FA_cout_236;
  (* register *) pwire FA_cout_237;
  (* register *) pwire FA_cout_238;
  (* register *) pwire FA_cout_239;
  (* register *) pwire FA_cout_240;
  (* register *) pwire FA_cout_241;
  (* register *) pwire FA_cout_242;
  (* register *) pwire FA_cout_243;
  (* register *) pwire FA_cout_244;
  (* register *) pwire FA_cout_245;
  (* register *) pwire FA_cout_246;
  (* register *) pwire FA_cout_247;
  (* register *) pwire FA_cout_248;
  (* register *) pwire FA_cout_249;
  (* register *) pwire FA_cout_250;
  (* register *) pwire FA_cout_251;
  (* register *) pwire FA_cout_252;
  (* register *) pwire FA_cout_253;
  (* register *) pwire FA_cout_254;
  (* register *) pwire FA_cout_255;
  (* register *) pwire FA_cout_256;
  (* register *) pwire FA_cout_257;
  (* register *) pwire FA_cout_258;
  (* register *) pwire FA_cout_259;
  (* register *) pwire FA_cout_260;
  (* register *) pwire FA_cout_261;
  (* register *) pwire FA_cout_262;
  (* register *) pwire FA_cout_263;
  (* register *) pwire FA_cout_264;
  (* register *) pwire FA_cout_265;
  (* register *) pwire FA_cout_266;
  (* register *) pwire FA_cout_267;
  (* register *) pwire FA_cout_268;
  (* register *) pwire FA_cout_269;
  (* register *) pwire FA_cout_270;
  (* register *) pwire FA_cout_271;
  (* register *) pwire FA_cout_272;
  (* register *) pwire FA_cout_273;
  (* register *) pwire FA_cout_274;
  (* register *) pwire FA_cout_275;
  (* register *) pwire FA_cout_276;
  (* register *) pwire FA_cout_277;
  (* register *) pwire FA_cout_278;
  (* register *) pwire FA_cout_279;
  (* register *) pwire FA_cout_280;
  (* register *) pwire FA_cout_281;
  (* register *) pwire FA_cout_282;
  (* register *) pwire FA_cout_283;
  (* register *) pwire FA_cout_284;
  (* register *) pwire FA_cout_285;
  (* register *) pwire FA_cout_286;
  (* register *) pwire FA_cout_287;
  (* register *) pwire FA_cout_288;
  (* register *) pwire FA_cout_289;
  (* register *) pwire FA_cout_290;
  (* register *) pwire FA_cout_291;
  (* register *) pwire FA_cout_292;
  (* register *) pwire FA_cout_293;
  (* register *) pwire FA_cout_294;
  (* register *) pwire FA_cout_295;
  (* register *) pwire FA_cout_296;
  (* register *) pwire FA_cout_297;
  (* register *) pwire FA_cout_298;
  (* register *) pwire FA_cout_299;
  (* register *) pwire FA_cout_300;
  (* register *) pwire FA_cout_301;
  (* register *) pwire FA_cout_302;
  (* register *) pwire FA_cout_303;
  (* register *) pwire FA_cout_304;
  (* register *) pwire FA_cout_305;
  (* register *) pwire FA_cout_306;
  (* register *) pwire FA_cout_307;
  (* register *) pwire FA_cout_308;
  (* register *) pwire FA_cout_309;
  (* register *) pwire FA_cout_310;
  (* register *) pwire FA_cout_311;
  (* register *) pwire FA_cout_312;
  (* register *) pwire FA_cout_313;
  (* register *) pwire FA_cout_314;
  (* register *) pwire FA_cout_315;
  (* register *) pwire FA_cout_316;
  (* register *) pwire FA_cout_317;
  (* register *) pwire FA_cout_318;
  (* register *) pwire FA_cout_319;
  (* register *) pwire FA_cout_320;
  (* register *) pwire FA_cout_321;
  (* register *) pwire FA_cout_322;
  (* register *) pwire FA_cout_323;
  (* register *) pwire FA_cout_324;
  (* register *) pwire FA_cout_325;
  (* register *) pwire FA_cout_326;
  (* register *) pwire FA_cout_327;
  (* register *) pwire FA_cout_328;
  (* register *) pwire FA_cout_329;
  (* register *) pwire FA_cout_330;
  (* register *) pwire FA_cout_331;
  (* register *) pwire FA_cout_332;
  (* register *) pwire FA_cout_333;
  (* register *) pwire FA_cout_334;
  (* register *) pwire FA_cout_335;
  (* register *) pwire FA_cout_336;
  (* register *) pwire FA_cout_337;
  (* register *) pwire FA_cout_338;
  (* register *) pwire FA_cout_339;
  (* register *) pwire FA_cout_340;
  (* register *) pwire FA_cout_341;
  (* register *) pwire FA_cout_342;
  (* register *) pwire FA_cout_343;
  (* register *) pwire FA_cout_344;
  (* register *) pwire FA_cout_345;
  (* register *) pwire FA_cout_346;
  (* register *) pwire FA_cout_347;
  (* register *) pwire FA_cout_348;
  (* register *) pwire FA_cout_349;
  (* register *) pwire FA_cout_350;
  (* register *) pwire FA_cout_351;
  (* register *) pwire FA_cout_352;
  (* register *) pwire FA_cout_353;
  (* register *) pwire FA_cout_354;
  (* register *) pwire FA_cout_355;
  (* register *) pwire FA_cout_356;
  (* register *) pwire FA_cout_357;
  (* register *) pwire FA_cout_358;
  (* register *) pwire FA_cout_359;
  (* register *) pwire FA_cout_360;
  (* register *) pwire FA_cout_361;
  (* register *) pwire FA_cout_362;
  (* register *) pwire FA_cout_363;
  (* register *) pwire FA_cout_364;
  (* register *) pwire FA_cout_365;
  (* register *) pwire FA_cout_366;
  (* register *) pwire FA_cout_367;
  (* register *) pwire FA_cout_368;
  (* register *) pwire FA_cout_369;
  (* register *) pwire FA_cout_370;
  (* register *) pwire FA_cout_371;
  (* register *) pwire FA_cout_372;
  (* register *) pwire FA_cout_373;
  (* register *) pwire FA_cout_374;
  (* register *) pwire FA_cout_375;
  (* register *) pwire FA_cout_376;
  (* register *) pwire FA_cout_377;
  (* register *) pwire FA_cout_378;
  (* register *) pwire FA_cout_379;
  (* register *) pwire FA_cout_380;
  (* register *) pwire FA_cout_381;
  (* register *) pwire FA_cout_382;
  (* register *) pwire FA_cout_383;
  (* register *) pwire FA_cout_384;
  (* register *) pwire FA_cout_385;
  (* register *) pwire FA_cout_386;
  (* register *) pwire FA_cout_387;
  (* register *) pwire FA_cout_388;
  (* register *) pwire FA_cout_389;
  (* register *) pwire FA_cout_390;
  (* register *) pwire FA_cout_391;
  (* register *) pwire FA_cout_392;
  (* register *) pwire FA_cout_393;
  (* register *) pwire FA_cout_394;
  (* register *) pwire FA_cout_395;
  (* register *) pwire FA_cout_396;
  (* register *) pwire FA_cout_397;
  (* register *) pwire FA_cout_398;
  (* register *) pwire FA_cout_399;
  (* register *) pwire FA_cout_400;
  (* register *) pwire FA_cout_401;
  (* register *) pwire FA_cout_402;
  (* register *) pwire FA_cout_403;
  (* register *) pwire FA_cout_404;
  (* register *) pwire FA_cout_405;
  (* register *) pwire FA_cout_406;
  (* register *) pwire FA_cout_407;
  (* register *) pwire FA_cout_408;
  (* register *) pwire FA_cout_409;
  (* register *) pwire FA_cout_410;
  (* register *) pwire FA_cout_411;
  (* register *) pwire FA_cout_412;
  (* register *) pwire FA_cout_413;
  (* register *) pwire FA_cout_414;
  (* register *) pwire FA_cout_415;
  (* register *) pwire FA_cout_416;
  (* register *) pwire FA_cout_417;
  (* register *) pwire FA_cout_418;
  (* register *) pwire FA_cout_419;
  (* register *) pwire FA_cout_420;
  (* register *) pwire FA_cout_421;
  (* register *) pwire FA_cout_422;
  (* register *) pwire FA_cout_423;
  (* register *) pwire FA_cout_424;
  (* register *) pwire FA_cout_425;
  (* register *) pwire FA_cout_426;
  (* register *) pwire FA_cout_427;
  (* register *) pwire FA_cout_428;
  (* register *) pwire FA_cout_429;
  (* register *) pwire FA_cout_430;
  (* register *) pwire FA_cout_431;
  (* register *) pwire FA_cout_432;
  (* register *) pwire FA_cout_433;
  (* register *) pwire FA_cout_434;
  (* register *) pwire FA_cout_435;
  (* register *) pwire FA_cout_436;
  (* register *) pwire FA_cout_437;
  (* register *) pwire FA_cout_438;
  (* register *) pwire FA_cout_439;
  (* register *) pwire FA_cout_440;
  (* register *) pwire FA_cout_441;
  (* register *) pwire FA_cout_442;
  (* register *) pwire FA_cout_443;
  (* register *) pwire FA_cout_444;
  (* register *) pwire FA_cout_445;
  (* register *) pwire FA_cout_446;
  (* register *) pwire FA_cout_447;
  (* register *) pwire FA_cout_448;
  (* register *) pwire FA_cout_449;
  (* register *) pwire FA_cout_450;
  (* register *) pwire FA_cout_451;
  (* register *) pwire FA_cout_452;
  (* register *) pwire FA_cout_453;
  (* register *) pwire FA_cout_454;
  (* register *) pwire FA_cout_455;
  (* register *) pwire FA_cout_456;
  (* register *) pwire FA_cout_457;
  (* register *) pwire FA_cout_458;
  (* register *) pwire FA_cout_459;
  (* register *) pwire FA_cout_460;
  (* register *) pwire FA_cout_461;
  (* register *) pwire FA_cout_462;
  (* register *) pwire FA_cout_463;
  (* register *) pwire FA_cout_464;
  (* register *) pwire FA_cout_465;
  (* register *) pwire FA_cout_466;
  (* register *) pwire FA_cout_467;
  (* register *) pwire FA_cout_468;
  (* register *) pwire FA_cout_469;
  (* register *) pwire FA_cout_470;
  (* register *) pwire FA_cout_471;
  (* register *) pwire FA_cout_472;
  (* register *) pwire FA_cout_473;
  (* register *) pwire FA_cout_474;
  (* register *) pwire FA_cout_475;
  (* register *) pwire FA_cout_476;
  (* register *) pwire FA_cout_477;
  (* register *) pwire FA_cout_478;
  (* register *) pwire FA_cout_479;
  (* register *) pwire FA_cout_480;
  (* register *) pwire FA_cout_481;
  (* register *) pwire FA_cout_482;
  (* register *) pwire FA_cout_483;
  (* register *) pwire FA_cout_484;
  (* register *) pwire FA_cout_485;
  (* register *) pwire FA_cout_486;
  (* register *) pwire FA_cout_487;
  (* register *) pwire FA_cout_488;
  (* register *) pwire FA_cout_489;
  (* register *) pwire FA_cout_490;
  (* register *) pwire FA_cout_491;
  (* register *) pwire FA_cout_492;
  (* register *) pwire FA_cout_493;
  (* register *) pwire FA_cout_494;
  (* register *) pwire FA_cout_495;
  (* register *) pwire FA_cout_496;
  (* register *) pwire FA_cout_497;
  (* register *) pwire FA_cout_498;
  (* register *) pwire FA_cout_499;
  (* register *) pwire FA_cout_500;
  (* register *) pwire FA_cout_501;
  (* register *) pwire FA_cout_502;
  (* register *) pwire FA_cout_503;
  (* register *) pwire FA_cout_504;
  (* register *) pwire FA_cout_505;
  (* register *) pwire FA_cout_506;
  (* register *) pwire FA_cout_507;
  (* register *) pwire FA_cout_508;
  (* register *) pwire FA_cout_509;
  (* register *) pwire FA_cout_510;
  (* register *) pwire FA_cout_511;
  (* register *) pwire FA_cout_512;
  (* register *) pwire FA_cout_513;
  (* register *) pwire FA_cout_514;
  (* register *) pwire FA_cout_515;
  (* register *) pwire FA_cout_516;
  (* register *) pwire FA_cout_517;
  (* register *) pwire FA_cout_518;
  (* register *) pwire FA_cout_519;
  (* register *) pwire FA_cout_520;
  (* register *) pwire FA_cout_521;
  (* register *) pwire FA_cout_522;
  (* register *) pwire FA_cout_523;
  (* register *) pwire FA_cout_524;
  (* register *) pwire FA_cout_525;
  (* register *) pwire FA_cout_526;
  (* register *) pwire FA_cout_527;
  (* register *) pwire FA_cout_528;
  (* register *) pwire FA_cout_529;
  (* register *) pwire FA_cout_530;
  (* register *) pwire FA_cout_531;
  (* register *) pwire FA_cout_532;
  (* register *) pwire FA_cout_533;
  (* register *) pwire FA_cout_534;
  (* register *) pwire FA_cout_535;
  (* register *) pwire FA_cout_536;
  (* register *) pwire FA_cout_537;
  (* register *) pwire FA_cout_538;
  (* register *) pwire FA_cout_539;
  (* register *) pwire FA_cout_540;
  (* register *) pwire FA_cout_541;
  (* register *) pwire FA_cout_542;
  (* register *) pwire FA_cout_543;
  (* register *) pwire FA_cout_544;
  (* register *) pwire FA_cout_545;
  (* register *) pwire FA_cout_546;
  (* register *) pwire FA_cout_547;
  (* register *) pwire FA_cout_548;
  (* register *) pwire FA_cout_549;
  (* register *) pwire FA_cout_550;
  (* register *) pwire FA_cout_551;
  (* register *) pwire FA_cout_552;
  (* register *) pwire FA_cout_553;
  (* register *) pwire FA_cout_554;
  (* register *) pwire FA_cout_555;
  (* register *) pwire FA_cout_556;
  (* register *) pwire FA_cout_557;
  (* register *) pwire FA_cout_558;
  (* register *) pwire FA_cout_559;
  (* register *) pwire FA_cout_560;
  (* register *) pwire FA_cout_561;
  (* register *) pwire FA_cout_562;
  (* register *) pwire FA_cout_563;
  (* register *) pwire FA_cout_564;
  (* register *) pwire FA_cout_565;
  (* register *) pwire FA_cout_566;
  (* register *) pwire FA_cout_567;
  (* register *) pwire FA_cout_568;
  (* register *) pwire FA_cout_569;
  (* register *) pwire FA_cout_570;
  (* register *) pwire FA_cout_571;
  (* register *) pwire FA_cout_572;
  (* register *) pwire FA_cout_573;
  (* register *) pwire FA_cout_574;
  (* register *) pwire FA_cout_575;
  (* register *) pwire FA_cout_576;
  (* register *) pwire FA_cout_577;
  (* register *) pwire FA_cout_578;
  (* register *) pwire FA_cout_579;
  (* register *) pwire FA_cout_580;
  (* register *) pwire FA_cout_581;
  (* register *) pwire FA_cout_582;
  (* register *) pwire FA_cout_583;
  (* register *) pwire FA_cout_584;
  (* register *) pwire FA_cout_585;
  (* register *) pwire FA_cout_586;
  (* register *) pwire FA_cout_587;
  (* register *) pwire FA_cout_588;
  (* register *) pwire FA_cout_589;
  (* register *) pwire FA_cout_590;
  (* register *) pwire FA_cout_591;
  (* register *) pwire FA_cout_592;
  (* register *) pwire FA_cout_593;
  (* register *) pwire FA_cout_594;
  (* register *) pwire FA_cout_595;
  (* register *) pwire FA_cout_596;
  (* register *) pwire FA_cout_597;
  (* register *) pwire FA_cout_598;
  (* register *) pwire FA_cout_599;
  (* register *) pwire FA_cout_600;
  (* register *) pwire FA_cout_601;
  (* register *) pwire FA_cout_602;
  (* register *) pwire FA_cout_603;
  (* register *) pwire FA_cout_604;
  (* register *) pwire FA_cout_605;
  (* register *) pwire FA_cout_606;
  (* register *) pwire FA_cout_607;
  (* register *) pwire FA_cout_608;
  (* register *) pwire FA_cout_609;
  (* register *) pwire FA_cout_610;
  (* register *) pwire FA_cout_611;
  (* register *) pwire FA_cout_612;
  (* register *) pwire FA_cout_613;
  (* register *) pwire FA_cout_614;
  (* register *) pwire FA_cout_615;
  (* register *) pwire FA_cout_616;
  (* register *) pwire FA_cout_617;
  (* register *) pwire FA_cout_618;
  (* register *) pwire FA_cout_619;
  (* register *) pwire FA_cout_620;
  (* register *) pwire FA_cout_621;
  (* register *) pwire FA_cout_622;
  (* register *) pwire FA_cout_623;
  (* register *) pwire FA_cout_624;
  (* register *) pwire FA_cout_625;
  (* register *) pwire FA_cout_626;
  (* register *) pwire FA_cout_627;
  (* register *) pwire FA_cout_628;
  (* register *) pwire FA_cout_629;
  (* register *) pwire FA_cout_630;
  (* register *) pwire FA_cout_631;
  (* register *) pwire FA_cout_632;
  (* register *) pwire FA_cout_633;
  (* register *) pwire FA_cout_634;
  (* register *) pwire FA_cout_635;
  (* register *) pwire FA_cout_636;
  (* register *) pwire FA_cout_637;
  (* register *) pwire FA_cout_638;
  (* register *) pwire FA_cout_639;
  (* register *) pwire FA_cout_640;
  (* register *) pwire FA_cout_641;
  (* register *) pwire FA_cout_642;
  (* register *) pwire FA_cout_643;
  (* register *) pwire FA_cout_644;
  (* register *) pwire FA_cout_645;
  (* register *) pwire FA_cout_646;
  (* register *) pwire FA_cout_647;
  (* register *) pwire FA_cout_648;
  (* register *) pwire FA_cout_649;
  (* register *) pwire FA_cout_650;
  (* register *) pwire FA_cout_651;
  (* register *) pwire FA_cout_652;
  (* register *) pwire FA_cout_653;
  (* register *) pwire FA_cout_654;
  (* register *) pwire FA_cout_655;
  (* register *) pwire FA_cout_656;
  (* register *) pwire FA_cout_657;
  (* register *) pwire FA_cout_658;
  (* register *) pwire FA_cout_659;
  (* register *) pwire FA_cout_660;
  (* register *) pwire FA_cout_661;
  (* register *) pwire FA_cout_662;
  (* register *) pwire FA_cout_663;
  (* register *) pwire FA_cout_664;
  (* register *) pwire FA_cout_665;
  (* register *) pwire FA_cout_666;
  (* register *) pwire FA_cout_667;
  (* register *) pwire FA_cout_668;
  (* register *) pwire FA_cout_669;
  (* register *) pwire FA_cout_670;
  (* register *) pwire FA_cout_671;
  (* register *) pwire FA_cout_672;
  (* register *) pwire FA_cout_673;
  (* register *) pwire FA_cout_674;
  (* register *) pwire FA_cout_675;
  (* register *) pwire FA_cout_676;
  (* register *) pwire FA_cout_677;
  (* register *) pwire FA_cout_678;
  (* register *) pwire FA_cout_679;
  (* register *) pwire FA_cout_680;
  (* register *) pwire FA_cout_681;
  (* register *) pwire FA_cout_682;
  (* register *) pwire FA_cout_683;
  (* register *) pwire FA_cout_684;
  (* register *) pwire FA_cout_685;
  (* register *) pwire FA_cout_686;
  (* register *) pwire FA_cout_687;
  (* register *) pwire FA_cout_688;
  (* register *) pwire FA_cout_689;
  (* register *) pwire FA_cout_690;
  (* register *) pwire FA_cout_691;
  (* register *) pwire FA_cout_692;
  (* register *) pwire FA_cout_693;
  (* register *) pwire FA_cout_694;
  (* register *) pwire FA_cout_695;
  (* register *) pwire FA_cout_696;
  (* register *) pwire FA_cout_697;
  (* register *) pwire FA_cout_698;
  (* register *) pwire FA_cout_699;
  (* register *) pwire FA_cout_700;
  (* register *) pwire FA_cout_701;
  (* register *) pwire FA_cout_702;
  (* register *) pwire FA_cout_703;
  (* register *) pwire FA_cout_704;
  (* register *) pwire FA_cout_705;
  (* register *) pwire FA_cout_706;
  (* register *) pwire FA_cout_707;
  (* register *) pwire FA_cout_708;
  (* register *) pwire FA_cout_709;
  (* register *) pwire FA_cout_710;
  (* register *) pwire FA_cout_711;
  (* register *) pwire FA_cout_712;
  (* register *) pwire FA_cout_713;
  (* register *) pwire FA_cout_714;
  (* register *) pwire FA_cout_715;
  (* register *) pwire FA_cout_716;
  (* register *) pwire FA_cout_717;
  (* register *) pwire FA_cout_718;
  (* register *) pwire FA_cout_719;
  (* register *) pwire FA_cout_720;
  (* register *) pwire FA_cout_721;
  (* register *) pwire FA_cout_722;
  (* register *) pwire FA_cout_723;
  (* register *) pwire FA_cout_724;
  (* register *) pwire FA_cout_725;
  (* register *) pwire FA_cout_726;
  (* register *) pwire FA_cout_727;
  (* register *) pwire FA_cout_728;
  (* register *) pwire FA_cout_729;
  (* register *) pwire FA_cout_730;
  (* register *) pwire FA_cout_731;
  (* register *) pwire FA_cout_732;
  (* register *) pwire FA_cout_733;
  (* register *) pwire FA_cout_734;
  (* register *) pwire FA_cout_735;
  (* register *) pwire FA_cout_736;
  (* register *) pwire FA_cout_737;
  (* register *) pwire FA_cout_738;
  (* register *) pwire FA_cout_739;
  (* register *) pwire FA_cout_740;
  (* register *) pwire FA_cout_741;
  (* register *) pwire FA_cout_742;
  (* register *) pwire FA_cout_743;
  (* register *) pwire FA_cout_744;
  (* register *) pwire FA_cout_745;
  (* register *) pwire FA_cout_746;
  (* register *) pwire FA_cout_747;
  (* register *) pwire FA_cout_748;
  (* register *) pwire FA_cout_749;
  (* register *) pwire FA_cout_750;
  (* register *) pwire FA_cout_751;
  (* register *) pwire FA_cout_752;
  (* register *) pwire FA_cout_753;
  (* register *) pwire FA_cout_754;
  (* register *) pwire FA_cout_755;
  (* register *) pwire FA_cout_756;
  (* register *) pwire FA_cout_757;
  (* register *) pwire FA_cout_758;
  (* register *) pwire FA_cout_759;
  (* register *) pwire FA_cout_760;
  (* register *) pwire FA_cout_761;
  (* register *) pwire FA_cout_762;
  (* register *) pwire FA_cout_763;
  (* register *) pwire FA_cout_764;
  (* register *) pwire FA_cout_765;
  (* register *) pwire FA_cout_766;
  (* register *) pwire FA_cout_767;
  (* register *) pwire FA_cout_768;
  (* register *) pwire FA_cout_769;
  (* register *) pwire FA_cout_770;
  (* register *) pwire FA_cout_771;
  (* register *) pwire FA_cout_772;
  (* register *) pwire FA_cout_773;
  (* register *) pwire FA_cout_774;
  (* register *) pwire FA_cout_775;
  (* register *) pwire FA_cout_776;
  (* register *) pwire FA_cout_777;
  (* register *) pwire FA_cout_778;
  (* register *) pwire FA_cout_779;
  (* register *) pwire FA_cout_780;
  (* register *) pwire FA_cout_781;
  (* register *) pwire FA_cout_782;
  (* register *) pwire FA_cout_783;
  (* register *) pwire FA_cout_784;
  (* register *) pwire FA_cout_785;
  (* register *) pwire FA_cout_786;
  (* register *) pwire FA_cout_787;
  (* register *) pwire FA_cout_788;
  (* register *) pwire FA_cout_789;
  (* register *) pwire FA_cout_790;
  (* register *) pwire FA_cout_791;
  (* register *) pwire FA_cout_792;
  (* register *) pwire FA_cout_793;
  (* register *) pwire FA_cout_794;
  (* register *) pwire FA_cout_795;
  (* register *) pwire FA_cout_796;
  (* register *) pwire FA_cout_797;
  (* register *) pwire FA_cout_798;
  (* register *) pwire FA_cout_799;
  (* register *) pwire FA_cout_800;
  (* register *) pwire FA_cout_801;
  (* register *) pwire FA_cout_802;
  (* register *) pwire FA_cout_803;
  (* register *) pwire FA_cout_804;
  (* register *) pwire FA_cout_805;
  (* register *) pwire FA_cout_806;
  (* register *) pwire FA_cout_807;
  (* register *) pwire FA_cout_808;
  (* register *) pwire FA_cout_809;
  (* register *) pwire FA_cout_810;
  (* register *) pwire FA_cout_811;
  (* register *) pwire FA_cout_812;
  (* register *) pwire FA_cout_813;
  (* register *) pwire FA_cout_814;
  (* register *) pwire FA_cout_815;
  (* register *) pwire FA_cout_816;
  (* register *) pwire FA_cout_817;
  (* register *) pwire FA_cout_818;
  (* register *) pwire FA_cout_819;
  (* register *) pwire FA_cout_820;
  (* register *) pwire FA_cout_821;
  (* register *) pwire FA_cout_822;
  (* register *) pwire FA_cout_823;
  (* register *) pwire FA_cout_824;
  (* register *) pwire FA_cout_825;
  (* register *) pwire FA_cout_826;
  (* register *) pwire FA_cout_827;
  (* register *) pwire FA_cout_828;
  (* register *) pwire FA_cout_829;
  (* register *) pwire FA_cout_830;
  (* register *) pwire FA_cout_831;
  (* register *) pwire FA_cout_832;
  (* register *) pwire FA_cout_833;
  (* register *) pwire FA_cout_834;
  (* register *) pwire FA_cout_835;
  (* register *) pwire FA_cout_836;
  (* register *) pwire FA_cout_837;
  (* register *) pwire FA_cout_838;
  (* register *) pwire FA_cout_839;
  (* register *) pwire FA_cout_840;
  (* register *) pwire FA_cout_841;
  (* register *) pwire FA_cout_842;
  (* register *) pwire FA_cout_843;
  (* register *) pwire FA_cout_844;
  (* register *) pwire FA_cout_845;
  (* register *) pwire FA_cout_846;
  (* register *) pwire FA_cout_847;
  (* register *) pwire FA_cout_848;
  (* register *) pwire FA_cout_849;
  (* register *) pwire FA_cout_850;
  (* register *) pwire FA_cout_851;
  (* register *) pwire FA_cout_852;
  (* register *) pwire FA_cout_853;
  (* register *) pwire FA_cout_854;
  (* register *) pwire FA_cout_855;
  (* register *) pwire FA_cout_856;
  (* register *) pwire FA_cout_857;
  (* register *) pwire FA_cout_858;
  (* register *) pwire FA_cout_859;
  (* register *) pwire FA_cout_860;
  (* register *) pwire FA_cout_861;
  (* register *) pwire FA_cout_862;
  (* register *) pwire FA_cout_863;
  (* register *) pwire FA_cout_864;
  (* register *) pwire FA_cout_865;
  (* register *) pwire FA_cout_866;
  (* register *) pwire FA_cout_867;
  (* register *) pwire FA_cout_868;
  (* register *) pwire FA_cout_869;
  (* register *) pwire FA_cout_870;
  (* register *) pwire FA_cout_871;
  (* register *) pwire FA_cout_872;
  (* register *) pwire FA_cout_873;
  (* register *) pwire FA_cout_874;
  (* register *) pwire FA_cout_875;
  (* register *) pwire FA_cout_876;
  (* register *) pwire FA_cout_877;
  (* register *) pwire FA_cout_878;
  (* register *) pwire FA_cout_879;
  (* register *) pwire FA_cout_880;
  (* register *) pwire FA_cout_881;
  (* register *) pwire FA_cout_882;
  (* register *) pwire FA_cout_883;
  (* register *) pwire FA_cout_884;
  (* register *) pwire FA_cout_885;
  (* register *) pwire FA_cout_886;
  (* register *) pwire FA_cout_887;
  (* register *) pwire FA_cout_888;
  (* register *) pwire FA_cout_889;
  (* register *) pwire FA_cout_890;
  (* register *) pwire FA_cout_891;
  (* register *) pwire FA_cout_892;
  (* register *) pwire FA_cout_893;
  (* register *) pwire FA_cout_894;
  (* register *) pwire FA_cout_895;
  (* register *) pwire FA_cout_896;
  (* register *) pwire FA_cout_897;
  (* register *) pwire FA_cout_898;
  (* register *) pwire FA_cout_899;
  (* register *) pwire FA_cout_900;
  (* register *) pwire FA_cout_901;
  (* register *) pwire FA_cout_902;
  (* register *) pwire FA_cout_903;
  (* register *) pwire FA_cout_904;
  (* register *) pwire FA_cout_905;
  (* register *) pwire FA_cout_906;
  (* register *) pwire FA_cout_907;
  (* register *) pwire FA_cout_908;
  (* register *) pwire FA_cout_909;
  (* register *) pwire FA_cout_910;
  (* register *) pwire FA_cout_911;
  (* register *) pwire FA_cout_912;
  (* register *) pwire FA_cout_913;
  (* register *) pwire FA_cout_914;
  (* register *) pwire FA_cout_915;
  (* register *) pwire FA_cout_916;
  (* register *) pwire FA_cout_917;
  (* register *) pwire FA_cout_918;
  (* register *) pwire FA_cout_919;
  (* register *) pwire FA_cout_920;
  (* register *) pwire FA_cout_921;
  (* register *) pwire FA_cout_922;
  (* register *) pwire FA_cout_923;
  (* register *) pwire FA_cout_924;
  (* register *) pwire FA_cout_925;
  (* register *) pwire FA_cout_926;
  (* register *) pwire FA_cout_927;
  (* register *) pwire FA_cout_928;
  (* register *) pwire FA_cout_929;
  (* register *) pwire FA_cout_930;
  (* register *) pwire FA_cout_931;
  (* register *) pwire FA_cout_932;
  (* register *) pwire FA_cout_933;
  (* register *) pwire FA_cout_934;
  (* register *) pwire FA_cout_935;
  (* register *) pwire FA_cout_936;
  (* register *) pwire FA_cout_937;
  (* register *) pwire FA_cout_938;
  (* register *) pwire FA_cout_939;
  (* register *) pwire FA_cout_940;
  (* register *) pwire FA_cout_941;
  (* register *) pwire FA_cout_942;
  (* register *) pwire FA_cout_943;
  (* register *) pwire FA_cout_944;
  (* register *) pwire FA_cout_945;
  (* register *) pwire FA_cout_946;
  (* register *) pwire FA_cout_947;
  (* register *) pwire FA_cout_948;
  (* register *) pwire FA_cout_949;
  (* register *) pwire FA_cout_950;
  (* register *) pwire FA_cout_951;
  (* register *) pwire FA_cout_952;
  (* register *) pwire FA_cout_953;
  (* register *) pwire FA_cout_954;
  (* register *) pwire FA_cout_955;
  (* register *) pwire FA_cout_956;
  (* register *) pwire FA_cout_957;
  (* register *) pwire FA_cout_958;
  (* register *) pwire FA_cout_959;
  (* register *) pwire FA_cout_960;
  (* register *) pwire FA_cout_961;
  (* register *) pwire FA_cout_962;
  (* register *) pwire FA_cout_963;
  (* register *) pwire FA_cout_964;
  (* register *) pwire FA_cout_965;
  (* register *) pwire FA_cout_966;
  (* register *) pwire FA_cout_967;
  (* register *) pwire FA_cout_968;
  (* register *) pwire FA_cout_969;
  (* register *) pwire FA_cout_970;
  (* register *) pwire FA_cout_971;
  (* register *) pwire FA_cout_972;
  (* register *) pwire FA_cout_973;
  (* register *) pwire FA_cout_974;
  (* register *) pwire FA_cout_975;
  (* register *) pwire FA_cout_976;
  (* register *) pwire FA_cout_977;
  (* register *) pwire FA_cout_978;
  (* register *) pwire FA_cout_979;
  (* register *) pwire FA_cout_980;
  (* register *) pwire FA_cout_981;
  (* register *) pwire FA_cout_982;
  (* register *) pwire FA_cout_983;
  (* register *) pwire FA_cout_984;
  (* register *) pwire FA_cout_985;
  (* register *) pwire FA_cout_986;
  (* register *) pwire FA_cout_987;
  (* register *) pwire FA_cout_988;
  (* register *) pwire FA_cout_989;
  (* register *) pwire FA_cout_990;
  (* register *) pwire FA_cout_991;
  (* register *) pwire FA_cout_992;
  (* register *) pwire FA_cout_993;
  (* register *) pwire FA_cout_994;
  (* register *) pwire FA_cout_995;
  (* register *) pwire FA_cout_996;
  (* register *) pwire FA_cout_997;
  (* register *) pwire FA_cout_998;
  (* register *) pwire FA_cout_999;
  (* register *) pwire FA_cout_1000;
  (* register *) pwire FA_cout_1001;
  (* register *) pwire FA_cout_1002;
  (* register *) pwire FA_cout_1003;
  (* register *) pwire FA_cout_1004;
  (* register *) pwire FA_cout_1005;
  (* register *) pwire FA_cout_1006;
  (* register *) pwire FA_cout_1007;
  (* register *) pwire FA_cout_1008;
  (* register *) pwire FA_cout_1009;
  (* register *) pwire FA_cout_1010;
  (* register *) pwire FA_cout_1011;
  (* register *) pwire FA_cout_1012;
  (* register *) pwire FA_cout_1013;
  (* register *) pwire FA_cout_1014;
  (* register *) pwire FA_cout_1015;
  (* register *) pwire FA_cout_1016;
  (* register *) pwire FA_cout_1017;
  (* register *) pwire FA_cout_1018;
  (* register *) pwire FA_cout_1019;
  (* register *) pwire FA_cout_1020;
  (* register *) pwire FA_cout_1021;
  (* register *) pwire FA_cout_1022;
  (* register *) pwire FA_cout_1023;
  (* register *) pwire FA_cout_1024;
  (* register *) pwire FA_cout_1025;
  (* register *) pwire FA_cout_1026;
  (* register *) pwire FA_cout_1027;
  (* register *) pwire FA_cout_1028;
  (* register *) pwire FA_cout_1029;
  (* register *) pwire FA_cout_1030;
  (* register *) pwire FA_cout_1031;
  (* register *) pwire FA_cout_1032;
  (* register *) pwire FA_cout_1033;
  (* register *) pwire FA_cout_1034;
  (* register *) pwire FA_cout_1035;
  (* register *) pwire FA_cout_1036;
  (* register *) pwire FA_cout_1037;
  (* register *) pwire FA_cout_1038;
  (* register *) pwire FA_cout_1039;
  (* register *) pwire FA_cout_1040;
  (* register *) pwire FA_cout_1041;
  (* register *) pwire FA_cout_1042;
  (* register *) pwire FA_cout_1043;
  (* register *) pwire FA_cout_1044;
  (* register *) pwire FA_cout_1045;
  (* register *) pwire FA_cout_1046;
  (* register *) pwire FA_cout_1047;
  (* register *) pwire FA_cout_1048;
  (* register *) pwire FA_cout_1049;
  (* register *) pwire FA_cout_1050;
  (* register *) pwire FA_cout_1051;
  (* register *) pwire FA_cout_1052;
  (* register *) pwire FA_cout_1053;
  (* register *) pwire FA_cout_1054;
  (* register *) pwire FA_cout_1055;
  (* register *) pwire FA_cout_1056;
  (* register *) pwire FA_cout_1057;
  (* register *) pwire FA_cout_1058;
  (* register *) pwire FA_cout_1059;
  (* register *) pwire FA_cout_1060;
  (* register *) pwire FA_cout_1061;
  (* register *) pwire FA_cout_1062;
  (* register *) pwire FA_cout_1063;
  (* register *) pwire FA_cout_1064;
  (* register *) pwire FA_cout_1065;
  (* register *) pwire FA_cout_1066;
  (* register *) pwire FA_cout_1067;
  (* register *) pwire FA_cout_1068;
  (* register *) pwire FA_cout_1069;
  (* register *) pwire FA_cout_1070;
  (* register *) pwire FA_cout_1071;
  (* register *) pwire FA_cout_1072;
  (* register *) pwire FA_cout_1073;
  (* register *) pwire FA_cout_1074;
  (* register *) pwire FA_cout_1075;
  (* register *) pwire FA_cout_1076;
  (* register *) pwire FA_cout_1077;
  (* register *) pwire FA_cout_1078;
  (* register *) pwire FA_cout_1079;
  (* register *) pwire FA_cout_1080;
  (* register *) pwire FA_cout_1081;
  (* register *) pwire FA_cout_1082;
  (* register *) pwire FA_cout_1083;
  (* register *) pwire FA_cout_1084;
  (* register *) pwire FA_cout_1085;
  (* register *) pwire FA_cout_1086;
  (* register *) pwire FA_cout_1087;
  (* register *) pwire FA_cout_1088;
  (* register *) pwire FA_cout_1089;
  (* register *) pwire FA_cout_1090;
  (* register *) pwire FA_cout_1091;
  (* register *) pwire FA_cout_1092;
  (* register *) pwire FA_cout_1093;
  (* register *) pwire FA_cout_1094;
  (* register *) pwire FA_cout_1095;
  (* register *) pwire FA_cout_1096;
  (* register *) pwire FA_cout_1097;
  (* register *) pwire FA_cout_1098;
  (* register *) pwire FA_cout_1099;
  (* register *) pwire FA_cout_1100;
  (* register *) pwire FA_cout_1101;
  (* register *) pwire FA_cout_1102;
  (* register *) pwire FA_cout_1103;
  (* register *) pwire FA_cout_1104;
  (* register *) pwire FA_cout_1105;
  (* register *) pwire FA_cout_1106;
  (* register *) pwire FA_cout_1107;
  (* register *) pwire FA_cout_1108;
  (* register *) pwire FA_cout_1109;
  (* register *) pwire FA_cout_1110;
  (* register *) pwire FA_cout_1111;
  (* register *) pwire FA_cout_1112;
  (* register *) pwire FA_cout_1113;
  (* register *) pwire FA_cout_1114;
  (* register *) pwire FA_cout_1115;
  (* register *) pwire FA_cout_1116;
  (* register *) pwire FA_cout_1117;
  (* register *) pwire FA_cout_1118;
  (* register *) pwire FA_cout_1119;
  (* register *) pwire FA_cout_1120;
  (* register *) pwire FA_cout_1121;
  (* register *) pwire FA_cout_1122;
  (* register *) pwire FA_cout_1123;
  (* register *) pwire FA_cout_1124;
  (* register *) pwire FA_cout_1125;
  (* register *) pwire FA_cout_1126;
  (* register *) pwire FA_cout_1127;
  (* register *) pwire FA_cout_1128;
  (* register *) pwire FA_cout_1129;
  (* register *) pwire FA_cout_1130;
  (* register *) pwire FA_cout_1131;
  (* register *) pwire FA_cout_1132;
  (* register *) pwire FA_cout_1133;
  (* register *) pwire FA_cout_1134;
  (* register *) pwire FA_cout_1135;
  (* register *) pwire FA_cout_1136;
  (* register *) pwire FA_cout_1137;
  (* register *) pwire FA_cout_1138;
  (* register *) pwire FA_cout_1139;
  (* register *) pwire FA_cout_1140;
  (* register *) pwire FA_cout_1141;
  (* register *) pwire FA_cout_1142;
  (* register *) pwire FA_cout_1143;
  (* register *) pwire FA_cout_1144;
  (* register *) pwire FA_cout_1145;
  (* register *) pwire FA_cout_1146;
  (* register *) pwire FA_cout_1147;
  (* register *) pwire FA_cout_1148;
  (* register *) pwire FA_cout_1149;
  (* register *) pwire FA_cout_1150;
  (* register *) pwire FA_cout_1151;
  (* register *) pwire FA_cout_1152;
  (* register *) pwire FA_cout_1153;
  (* register *) pwire FA_cout_1154;
  (* register *) pwire FA_cout_1155;
  (* register *) pwire FA_cout_1156;
  (* register *) pwire FA_cout_1157;
  (* register *) pwire FA_cout_1158;
  (* register *) pwire FA_cout_1159;
  (* register *) pwire FA_cout_1160;
  (* register *) pwire FA_cout_1161;
  (* register *) pwire FA_cout_1162;
  (* register *) pwire FA_cout_1163;
  (* register *) pwire FA_cout_1164;
  (* register *) pwire FA_cout_1165;
  (* register *) pwire FA_cout_1166;
  (* register *) pwire FA_cout_1167;
  (* register *) pwire FA_cout_1168;
  (* register *) pwire FA_cout_1169;
  (* register *) pwire FA_cout_1170;
  (* register *) pwire FA_cout_1171;
  (* register *) pwire FA_cout_1172;
  (* register *) pwire FA_cout_1173;
  (* register *) pwire FA_cout_1174;
  (* register *) pwire FA_cout_1175;
  (* register *) pwire FA_cout_1176;
  (* register *) pwire FA_cout_1177;
  (* register *) pwire FA_cout_1178;
  (* register *) pwire FA_cout_1179;
  (* register *) pwire FA_cout_1180;
  (* register *) pwire FA_cout_1181;
  (* register *) pwire FA_cout_1182;
  (* register *) pwire FA_cout_1183;
  (* register *) pwire FA_cout_1184;
  (* register *) pwire FA_cout_1185;
  (* register *) pwire FA_cout_1186;
  (* register *) pwire FA_cout_1187;
  (* register *) pwire FA_cout_1188;
  (* register *) pwire FA_cout_1189;
  (* register *) pwire FA_cout_1190;
  (* register *) pwire FA_cout_1191;
  (* register *) pwire FA_cout_1192;
  (* register *) pwire FA_cout_1193;
  (* register *) pwire FA_cout_1194;
  (* register *) pwire FA_cout_1195;
  (* register *) pwire FA_cout_1196;
  (* register *) pwire FA_cout_1197;
  (* register *) pwire FA_cout_1198;
  (* register *) pwire FA_cout_1199;
  (* register *) pwire FA_cout_1200;
  (* register *) pwire FA_cout_1201;
  (* register *) pwire FA_cout_1202;
  (* register *) pwire FA_cout_1203;
  (* register *) pwire FA_cout_1204;
  (* register *) pwire FA_cout_1205;
  (* register *) pwire FA_cout_1206;
  (* register *) pwire FA_cout_1207;
  (* register *) pwire FA_cout_1208;
  (* register *) pwire FA_cout_1209;
  (* register *) pwire FA_cout_1210;
  (* register *) pwire FA_cout_1211;
  (* register *) pwire FA_cout_1212;
  (* register *) pwire FA_cout_1213;
  (* register *) pwire FA_cout_1214;
  (* register *) pwire FA_cout_1215;
  (* register *) pwire FA_cout_1216;
  (* register *) pwire FA_cout_1217;
  (* register *) pwire FA_cout_1218;
  (* register *) pwire FA_cout_1219;
  (* register *) pwire FA_cout_1220;
  (* register *) pwire FA_cout_1221;
  (* register *) pwire FA_cout_1222;
  (* register *) pwire FA_cout_1223;
  (* register *) pwire FA_cout_1224;
  (* register *) pwire FA_cout_1225;
  (* register *) pwire FA_cout_1226;
  (* register *) pwire FA_cout_1227;
  (* register *) pwire FA_cout_1228;
  (* register *) pwire FA_cout_1229;
  (* register *) pwire FA_cout_1230;
  (* register *) pwire FA_cout_1231;
  (* register *) pwire FA_cout_1232;
  (* register *) pwire FA_cout_1233;
  (* register *) pwire FA_cout_1234;
  (* register *) pwire FA_cout_1235;
  (* register *) pwire FA_cout_1236;
  (* register *) pwire FA_cout_1237;
  (* register *) pwire FA_cout_1238;
  (* register *) pwire FA_cout_1239;
  (* register *) pwire FA_cout_1240;
  (* register *) pwire FA_cout_1241;
  (* register *) pwire FA_cout_1242;
  (* register *) pwire FA_cout_1243;
  (* register *) pwire FA_cout_1244;
  (* register *) pwire FA_cout_1245;
  (* register *) pwire FA_cout_1246;
  (* register *) pwire FA_cout_1247;
  (* register *) pwire FA_cout_1248;
  (* register *) pwire FA_cout_1249;
  (* register *) pwire FA_cout_1250;
  (* register *) pwire FA_cout_1251;
  (* register *) pwire FA_cout_1252;
  (* register *) pwire FA_cout_1253;
  (* register *) pwire FA_cout_1254;
  (* register *) pwire FA_cout_1255;
  (* register *) pwire FA_cout_1256;
  (* register *) pwire FA_cout_1257;
  (* register *) pwire FA_cout_1258;
  (* register *) pwire FA_cout_1259;
  (* register *) pwire FA_cout_1260;
  (* register *) pwire FA_cout_1261;
  (* register *) pwire FA_cout_1262;
  (* register *) pwire FA_cout_1263;
  (* register *) pwire FA_cout_1264;
  (* register *) pwire FA_cout_1265;
  (* register *) pwire FA_cout_1266;
  (* register *) pwire FA_cout_1267;
  (* register *) pwire FA_cout_1268;
  (* register *) pwire FA_cout_1269;
  (* register *) pwire FA_cout_1270;
  (* register *) pwire FA_cout_1271;
  (* register *) pwire FA_cout_1272;
  (* register *) pwire FA_cout_1273;
  (* register *) pwire FA_cout_1274;
  (* register *) pwire FA_cout_1275;
  (* register *) pwire FA_cout_1276;
  (* register *) pwire FA_cout_1277;
  (* register *) pwire FA_cout_1278;
  (* register *) pwire FA_cout_1279;
  (* register *) pwire FA_cout_1280;
  (* register *) pwire FA_cout_1281;
  (* register *) pwire FA_cout_1282;
  (* register *) pwire FA_cout_1283;
  (* register *) pwire FA_cout_1284;
  (* register *) pwire FA_cout_1285;
  (* register *) pwire FA_cout_1286;
  (* register *) pwire FA_cout_1287;
  (* register *) pwire FA_cout_1288;
  (* register *) pwire FA_cout_1289;
  (* register *) pwire FA_cout_1290;
  (* register *) pwire FA_cout_1291;
  (* register *) pwire FA_cout_1292;
  (* register *) pwire FA_cout_1293;
  (* register *) pwire FA_cout_1294;
  (* register *) pwire FA_cout_1295;
  (* register *) pwire FA_cout_1296;
  (* register *) pwire FA_cout_1297;
  (* register *) pwire FA_cout_1298;
  (* register *) pwire FA_cout_1299;
  (* register *) pwire FA_cout_1300;
  (* register *) pwire FA_cout_1301;
  (* register *) pwire FA_cout_1302;
  (* register *) pwire FA_cout_1303;
  (* register *) pwire FA_cout_1304;
  (* register *) pwire FA_cout_1305;
  (* register *) pwire FA_cout_1306;
  (* register *) pwire FA_cout_1307;
  (* register *) pwire FA_cout_1308;
  (* register *) pwire FA_cout_1309;
  (* register *) pwire FA_cout_1310;
  (* register *) pwire FA_cout_1311;
  (* register *) pwire FA_cout_1312;
  (* register *) pwire FA_cout_1313;
  (* register *) pwire FA_cout_1314;
  (* register *) pwire FA_cout_1315;
  (* register *) pwire FA_cout_1316;
  (* register *) pwire FA_cout_1317;
  (* register *) pwire FA_cout_1318;
  (* register *) pwire FA_cout_1319;
  (* register *) pwire FA_cout_1320;
  (* register *) pwire FA_cout_1321;
  (* register *) pwire FA_cout_1322;
  (* register *) pwire FA_cout_1323;
  (* register *) pwire FA_cout_1324;
  (* register *) pwire FA_cout_1325;
  (* register *) pwire FA_cout_1326;
  (* register *) pwire FA_cout_1327;
  (* register *) pwire FA_cout_1328;
  (* register *) pwire FA_cout_1329;
  (* register *) pwire FA_cout_1330;
  (* register *) pwire FA_cout_1331;
  (* register *) pwire FA_cout_1332;
  (* register *) pwire FA_cout_1333;
  (* register *) pwire FA_cout_1334;
  (* register *) pwire FA_cout_1335;
  (* register *) pwire FA_cout_1336;
  (* register *) pwire FA_cout_1337;
  (* register *) pwire FA_cout_1338;
  (* register *) pwire FA_cout_1339;
  (* register *) pwire FA_cout_1340;
  (* register *) pwire FA_cout_1341;
  (* register *) pwire FA_cout_1342;
  (* register *) pwire FA_cout_1343;
  (* register *) pwire FA_cout_1344;
  (* register *) pwire FA_cout_1345;
  (* register *) pwire FA_cout_1346;
  (* register *) pwire FA_cout_1347;
  (* register *) pwire FA_cout_1348;
  (* register *) pwire FA_cout_1349;
  (* register *) pwire FA_cout_1350;
  (* register *) pwire FA_cout_1351;
  (* register *) pwire FA_cout_1352;
  (* register *) pwire FA_cout_1353;
  (* register *) pwire FA_cout_1354;
  (* register *) pwire FA_cout_1355;
  (* register *) pwire FA_cout_1356;
  (* register *) pwire FA_cout_1357;
  (* register *) pwire FA_cout_1358;
  (* register *) pwire FA_cout_1359;
  (* register *) pwire FA_cout_1360;
  (* register *) pwire FA_cout_1361;
  (* register *) pwire FA_cout_1362;
  (* register *) pwire FA_cout_1363;
  (* register *) pwire FA_cout_1364;
  (* register *) pwire FA_cout_1365;
  (* register *) pwire FA_cout_1366;
  (* register *) pwire FA_cout_1367;
  (* register *) pwire FA_cout_1368;
  (* register *) pwire FA_cout_1369;
  (* register *) pwire FA_cout_1370;
  (* register *) pwire FA_cout_1371;
  (* register *) pwire FA_cout_1372;
  (* register *) pwire FA_cout_1373;
  (* register *) pwire FA_cout_1374;
  (* register *) pwire FA_cout_1375;
  (* register *) pwire FA_cout_1376;
  (* register *) pwire FA_cout_1377;
  (* register *) pwire FA_cout_1378;
  (* register *) pwire FA_cout_1379;
  (* register *) pwire FA_cout_1380;
  (* register *) pwire FA_cout_1381;
  (* register *) pwire FA_cout_1382;
  (* register *) pwire FA_cout_1383;
  (* register *) pwire FA_cout_1384;
  (* register *) pwire FA_cout_1385;
  (* register *) pwire FA_cout_1386;
  (* register *) pwire FA_cout_1387;
  (* register *) pwire FA_cout_1388;
  (* register *) pwire FA_cout_1389;
  (* register *) pwire FA_cout_1390;
  (* register *) pwire FA_cout_1391;
  (* register *) pwire FA_cout_1392;
  (* register *) pwire FA_cout_1393;
  (* register *) pwire FA_cout_1394;
  (* register *) pwire FA_cout_1395;
  (* register *) pwire FA_cout_1396;
  (* register *) pwire FA_cout_1397;
  (* register *) pwire FA_cout_1398;
  (* register *) pwire FA_cout_1399;
  (* register *) pwire FA_cout_1400;
  (* register *) pwire FA_cout_1401;
  (* register *) pwire FA_cout_1402;
  (* register *) pwire FA_cout_1403;
  (* register *) pwire FA_cout_1404;
  (* register *) pwire FA_cout_1405;
  (* register *) pwire FA_cout_1406;
  (* register *) pwire FA_cout_1407;
  (* register *) pwire FA_cout_1408;
  (* register *) pwire FA_cout_1409;
  (* register *) pwire FA_cout_1410;
  (* register *) pwire FA_cout_1411;
  (* register *) pwire FA_cout_1412;
  (* register *) pwire FA_cout_1413;
  (* register *) pwire FA_cout_1414;
  (* register *) pwire FA_cout_1415;
  (* register *) pwire FA_cout_1416;
  (* register *) pwire FA_cout_1417;
  (* register *) pwire FA_cout_1418;
  (* register *) pwire FA_cout_1419;
  (* register *) pwire FA_cout_1420;
  (* register *) pwire FA_cout_1421;
  (* register *) pwire FA_cout_1422;
  (* register *) pwire FA_cout_1423;
  (* register *) pwire FA_cout_1424;
  (* register *) pwire FA_cout_1425;
  (* register *) pwire FA_cout_1426;
  (* register *) pwire FA_cout_1427;
  (* register *) pwire FA_cout_1428;
  (* register *) pwire FA_cout_1429;
  (* register *) pwire FA_cout_1430;
  (* register *) pwire FA_cout_1431;
  (* register *) pwire FA_cout_1432;
  (* register *) pwire FA_cout_1433;
  (* register *) pwire FA_cout_1434;
  (* register *) pwire FA_cout_1435;
  (* register *) pwire FA_cout_1436;
  (* register *) pwire FA_cout_1437;
  (* register *) pwire FA_cout_1438;
  (* register *) pwire FA_cout_1439;
  (* register *) pwire FA_cout_1440;
  (* register *) pwire FA_cout_1441;
  (* register *) pwire FA_cout_1442;
  (* register *) pwire FA_cout_1443;
  (* register *) pwire FA_cout_1444;
  (* register *) pwire FA_cout_1445;
  (* register *) pwire FA_cout_1446;
  (* register *) pwire FA_cout_1447;
  (* register *) pwire FA_cout_1448;
  (* register *) pwire FA_cout_1449;
  (* register *) pwire FA_cout_1450;
  (* register *) pwire FA_cout_1451;
  (* register *) pwire FA_cout_1452;
  (* register *) pwire FA_cout_1453;
  (* register *) pwire FA_cout_1454;
  (* register *) pwire FA_cout_1455;
  (* register *) pwire FA_cout_1456;
  (* register *) pwire FA_cout_1457;
  (* register *) pwire FA_cout_1458;
  (* register *) pwire FA_cout_1459;
  (* register *) pwire FA_cout_1460;
  (* register *) pwire FA_cout_1461;
  (* register *) pwire FA_cout_1462;
  (* register *) pwire FA_cout_1463;
  (* register *) pwire FA_cout_1464;
  (* register *) pwire FA_cout_1465;
  (* register *) pwire FA_cout_1466;
  (* register *) pwire FA_cout_1467;
  (* register *) pwire FA_cout_1468;
  (* register *) pwire FA_cout_1469;
  (* register *) pwire FA_cout_1470;
  (* register *) pwire FA_cout_1471;
  (* register *) pwire FA_cout_1472;
  (* register *) pwire FA_cout_1473;
  (* register *) pwire FA_cout_1474;
  (* register *) pwire FA_cout_1475;
  (* register *) pwire FA_cout_1476;
  (* register *) pwire FA_cout_1477;
  (* register *) pwire FA_cout_1478;
  (* register *) pwire FA_cout_1479;
  (* register *) pwire FA_cout_1480;
  (* register *) pwire FA_cout_1481;
  (* register *) pwire FA_cout_1482;
  (* register *) pwire FA_cout_1483;
  (* register *) pwire FA_cout_1484;
  (* register *) pwire FA_cout_1485;
  (* register *) pwire FA_cout_1486;
  (* register *) pwire FA_cout_1487;
  (* register *) pwire FA_cout_1488;
  (* register *) pwire FA_cout_1489;
  (* register *) pwire FA_cout_1490;
  (* register *) pwire FA_cout_1491;
  (* register *) pwire FA_cout_1492;
  (* register *) pwire FA_cout_1493;
  (* register *) pwire FA_cout_1494;
  (* register *) pwire FA_cout_1495;
  (* register *) pwire FA_cout_1496;
  (* register *) pwire FA_cout_1497;
  (* register *) pwire FA_cout_1498;
  (* register *) pwire FA_cout_1499;
  (* register *) pwire FA_cout_1500;
  (* register *) pwire FA_cout_1501;
  (* register *) pwire FA_cout_1502;
  (* register *) pwire FA_cout_1503;
  (* register *) pwire FA_cout_1504;
  (* register *) pwire FA_cout_1505;
  (* register *) pwire FA_cout_1506;
  (* register *) pwire FA_cout_1507;
  (* register *) pwire FA_cout_1508;
  (* register *) pwire FA_cout_1509;
  (* register *) pwire FA_cout_1510;
  (* register *) pwire FA_cout_1511;
  (* register *) pwire FA_cout_1512;
  (* register *) pwire FA_cout_1513;
  (* register *) pwire FA_cout_1514;
  (* register *) pwire FA_cout_1515;
  (* register *) pwire FA_cout_1516;
  (* register *) pwire FA_cout_1517;
  (* register *) pwire FA_cout_1518;
  (* register *) pwire FA_cout_1519;
  (* register *) pwire FA_cout_1520;
  (* register *) pwire FA_cout_1521;
  (* register *) pwire FA_cout_1522;
  (* register *) pwire FA_cout_1523;
  (* register *) pwire FA_cout_1524;
  (* register *) pwire FA_cout_1525;
  (* register *) pwire FA_cout_1526;
  (* register *) pwire FA_cout_1527;
  (* register *) pwire FA_cout_1528;
  (* register *) pwire FA_cout_1529;
  (* register *) pwire FA_cout_1530;
  (* register *) pwire FA_cout_1531;
  (* register *) pwire FA_cout_1532;
  (* register *) pwire FA_cout_1533;
  (* register *) pwire FA_cout_1534;
  (* register *) pwire FA_cout_1535;
  (* register *) pwire FA_cout_1536;
  (* register *) pwire FA_cout_1537;
  (* register *) pwire FA_cout_1538;
  (* register *) pwire FA_cout_1539;
  (* register *) pwire FA_cout_1540;
  (* register *) pwire FA_cout_1541;
  (* register *) pwire FA_cout_1542;
  (* register *) pwire FA_cout_1543;
  (* register *) pwire FA_cout_1544;
  (* register *) pwire FA_cout_1545;
  (* register *) pwire FA_cout_1546;
  (* register *) pwire FA_cout_1547;
  (* register *) pwire FA_cout_1548;
  (* register *) pwire FA_cout_1549;
  (* register *) pwire FA_cout_1550;
  (* register *) pwire FA_cout_1551;
  (* register *) pwire FA_cout_1552;
  (* register *) pwire FA_cout_1553;
  (* register *) pwire FA_cout_1554;
  (* register *) pwire FA_cout_1555;
  (* register *) pwire FA_cout_1556;
  (* register *) pwire FA_cout_1557;
  (* register *) pwire FA_cout_1558;
  (* register *) pwire FA_cout_1559;
  (* register *) pwire FA_cout_1560;
  (* register *) pwire FA_cout_1561;
  (* register *) pwire FA_cout_1562;
  (* register *) pwire FA_cout_1563;
  (* register *) pwire FA_cout_1564;
  (* register *) pwire FA_cout_1565;
  (* register *) pwire FA_cout_1566;
  (* register *) pwire FA_cout_1567;
  (* register *) pwire FA_cout_1568;
  (* register *) pwire FA_cout_1569;
  (* register *) pwire FA_cout_1570;
  (* register *) pwire FA_cout_1571;
  (* register *) pwire FA_cout_1572;
  (* register *) pwire FA_cout_1573;
  (* register *) pwire FA_cout_1574;
  (* register *) pwire FA_cout_1575;
  (* register *) pwire FA_cout_1576;
  (* register *) pwire FA_cout_1577;
  (* register *) pwire FA_cout_1578;
  (* register *) pwire FA_cout_1579;
  (* register *) pwire FA_cout_1580;
  (* register *) pwire FA_cout_1581;
  (* register *) pwire FA_cout_1582;
  (* register *) pwire FA_cout_1583;
  (* register *) pwire FA_cout_1584;
  (* register *) pwire FA_cout_1585;
  (* register *) pwire FA_cout_1586;
  (* register *) pwire FA_cout_1587;
  (* register *) pwire FA_cout_1588;
  (* register *) pwire FA_cout_1589;
  (* register *) pwire FA_cout_1590;
  (* register *) pwire FA_cout_1591;
  (* register *) pwire FA_cout_1592;
  (* register *) pwire FA_cout_1593;
  (* register *) pwire FA_cout_1594;
  (* register *) pwire FA_cout_1595;
  (* register *) pwire FA_cout_1596;
  (* register *) pwire FA_cout_1597;
  (* register *) pwire FA_cout_1598;
  (* register *) pwire FA_cout_1599;
  (* register *) pwire FA_cout_1600;
  (* register *) pwire FA_cout_1601;
  (* register *) pwire FA_cout_1602;
  (* register *) pwire FA_cout_1603;
  (* register *) pwire FA_cout_1604;
  (* register *) pwire FA_cout_1605;
  (* register *) pwire FA_cout_1606;
  (* register *) pwire FA_cout_1607;
  (* register *) pwire FA_cout_1608;
  (* register *) pwire FA_cout_1609;
  (* register *) pwire FA_cout_1610;
  (* register *) pwire FA_cout_1611;
  (* register *) pwire FA_cout_1612;
  (* register *) pwire FA_cout_1613;
  (* register *) pwire FA_cout_1614;
  (* register *) pwire FA_cout_1615;
  (* register *) pwire FA_cout_1616;
  (* register *) pwire FA_cout_1617;
  (* register *) pwire FA_cout_1618;
  (* register *) pwire FA_cout_1619;
  (* register *) pwire FA_cout_1620;
  (* register *) pwire FA_cout_1621;
  (* register *) pwire FA_cout_1622;
  (* register *) pwire FA_cout_1623;
  (* register *) pwire FA_cout_1624;
  (* register *) pwire FA_cout_1625;
  (* register *) pwire FA_cout_1626;
  (* register *) pwire FA_cout_1627;
  (* register *) pwire FA_cout_1628;
  (* register *) pwire FA_cout_1629;
  (* register *) pwire FA_cout_1630;
  (* register *) pwire FA_cout_1631;
  (* register *) pwire FA_cout_1632;
  (* register *) pwire FA_cout_1633;
  (* register *) pwire FA_cout_1634;
  (* register *) pwire FA_cout_1635;
  (* register *) pwire FA_cout_1636;
  (* register *) pwire FA_cout_1637;
  (* register *) pwire FA_cout_1638;
  (* register *) pwire FA_cout_1639;
  (* register *) pwire FA_cout_1640;
  (* register *) pwire FA_cout_1641;
  (* register *) pwire FA_cout_1642;
  (* register *) pwire FA_cout_1643;
  (* register *) pwire FA_cout_1644;
  (* register *) pwire FA_cout_1645;
  (* register *) pwire FA_cout_1646;
  (* register *) pwire FA_cout_1647;
  (* register *) pwire FA_cout_1648;
  (* register *) pwire FA_cout_1649;
  (* register *) pwire FA_cout_1650;
  (* register *) pwire FA_cout_1651;
  (* register *) pwire FA_cout_1652;
  (* register *) pwire FA_cout_1653;
  (* register *) pwire FA_cout_1654;
  (* register *) pwire FA_cout_1655;
  (* register *) pwire FA_cout_1656;
  (* register *) pwire FA_cout_1657;
  (* register *) pwire FA_cout_1658;
  (* register *) pwire FA_cout_1659;
  (* register *) pwire FA_cout_1660;
  (* register *) pwire FA_cout_1661;
  (* register *) pwire FA_cout_1662;
  (* register *) pwire FA_cout_1663;
  (* register *) pwire FA_cout_1664;
  (* register *) pwire FA_cout_1665;
  (* register *) pwire FA_cout_1666;
  (* register *) pwire FA_cout_1667;
  (* register *) pwire FA_cout_1668;
  (* register *) pwire FA_cout_1669;
  (* register *) pwire FA_cout_1670;
  (* register *) pwire FA_cout_1671;
  (* register *) pwire FA_cout_1672;
  (* register *) pwire FA_cout_1673;
  (* register *) pwire FA_cout_1674;
  (* register *) pwire FA_cout_1675;
  (* register *) pwire FA_cout_1676;
  (* register *) pwire FA_cout_1677;
  (* register *) pwire FA_cout_1678;
  (* register *) pwire FA_cout_1679;
  (* register *) pwire FA_cout_1680;
  (* register *) pwire FA_cout_1681;
  (* register *) pwire FA_cout_1682;
  (* register *) pwire FA_cout_1683;
  (* register *) pwire FA_cout_1684;
  (* register *) pwire FA_cout_1685;
  (* register *) pwire FA_cout_1686;
  (* register *) pwire FA_cout_1687;
  (* register *) pwire FA_cout_1688;
  (* register *) pwire FA_cout_1689;
  (* register *) pwire FA_cout_1690;
  (* register *) pwire FA_cout_1691;
  (* register *) pwire FA_cout_1692;
  (* register *) pwire FA_cout_1693;
  (* register *) pwire FA_cout_1694;
  (* register *) pwire FA_cout_1695;
  (* register *) pwire FA_cout_1696;
  (* register *) pwire FA_cout_1697;
  (* register *) pwire FA_cout_1698;
  (* register *) pwire FA_cout_1699;
  (* register *) pwire FA_cout_1700;
  (* register *) pwire FA_cout_1701;
  (* register *) pwire FA_cout_1702;
  (* register *) pwire FA_cout_1703;
  (* register *) pwire FA_cout_1704;
  (* register *) pwire FA_cout_1705;
  (* register *) pwire FA_cout_1706;
  (* register *) pwire FA_cout_1707;
  (* register *) pwire FA_cout_1708;
  (* register *) pwire FA_cout_1709;
  (* register *) pwire FA_cout_1710;
  (* register *) pwire FA_cout_1711;
  (* register *) pwire FA_cout_1712;
  (* register *) pwire FA_cout_1713;
  (* register *) pwire FA_cout_1714;
  (* register *) pwire FA_cout_1715;
  (* register *) pwire FA_cout_1716;
  (* register *) pwire FA_cout_1717;
  (* register *) pwire FA_cout_1718;
  (* register *) pwire FA_cout_1719;
  (* register *) pwire FA_cout_1720;
  (* register *) pwire FA_cout_1721;
  (* register *) pwire FA_cout_1722;
  (* register *) pwire FA_cout_1723;
  (* register *) pwire FA_cout_1724;
  (* register *) pwire FA_cout_1725;
  (* register *) pwire FA_cout_1726;
  (* register *) pwire FA_cout_1727;
  (* register *) pwire FA_cout_1728;
  (* register *) pwire FA_cout_1729;
  (* register *) pwire FA_cout_1730;
  (* register *) pwire FA_cout_1731;
  (* register *) pwire FA_cout_1732;
  (* register *) pwire FA_cout_1733;
  (* register *) pwire FA_cout_1734;
  (* register *) pwire FA_cout_1735;
  (* register *) pwire FA_cout_1736;
  (* register *) pwire FA_cout_1737;
  (* register *) pwire FA_cout_1738;
  (* register *) pwire FA_cout_1739;
  (* register *) pwire FA_cout_1740;
  (* register *) pwire FA_cout_1741;
  (* register *) pwire FA_cout_1742;
  (* register *) pwire FA_cout_1743;
  (* register *) pwire FA_cout_1744;
  (* register *) pwire FA_cout_1745;
  (* register *) pwire FA_cout_1746;
  (* register *) pwire FA_cout_1747;
  (* register *) pwire FA_cout_1748;
  (* register *) pwire FA_cout_1749;
  (* register *) pwire FA_cout_1750;
  (* register *) pwire FA_cout_1751;
  (* register *) pwire FA_cout_1752;
  (* register *) pwire FA_cout_1753;
  (* register *) pwire FA_cout_1754;
  (* register *) pwire FA_cout_1755;
  (* register *) pwire FA_cout_1756;
  (* register *) pwire FA_cout_1757;
  (* register *) pwire FA_cout_1758;
  (* register *) pwire FA_cout_1759;
  (* register *) pwire FA_cout_1760;
  (* register *) pwire FA_cout_1761;
  (* register *) pwire FA_cout_1762;
  (* register *) pwire FA_cout_1763;
  (* register *) pwire FA_cout_1764;
  (* register *) pwire FA_cout_1765;
  (* register *) pwire FA_cout_1766;
  (* register *) pwire FA_cout_1767;
  (* register *) pwire FA_cout_1768;
  (* register *) pwire FA_cout_1769;
  (* register *) pwire FA_cout_1770;
  (* register *) pwire FA_cout_1771;
  (* register *) pwire FA_cout_1772;
  (* register *) pwire FA_cout_1773;
  (* register *) pwire FA_cout_1774;
  (* register *) pwire FA_cout_1775;
  (* register *) pwire FA_cout_1776;
  (* register *) pwire FA_cout_1777;
  (* register *) pwire FA_cout_1778;
  (* register *) pwire FA_cout_1779;
  (* register *) pwire FA_cout_1780;
  (* register *) pwire FA_cout_1781;
  (* register *) pwire FA_cout_1782;
  (* register *) pwire FA_cout_1783;
  (* register *) pwire FA_cout_1784;
  (* register *) pwire FA_cout_1785;
  (* register *) pwire FA_cout_1786;
  (* register *) pwire FA_cout_1787;
  (* register *) pwire FA_cout_1788;
  (* register *) pwire FA_cout_1789;
  (* register *) pwire FA_cout_1790;
  (* register *) pwire FA_cout_1791;
  (* register *) pwire FA_cout_1792;
  (* register *) pwire FA_cout_1793;
  (* register *) pwire FA_cout_1794;
  (* register *) pwire FA_cout_1795;
  (* register *) pwire FA_cout_1796;
  (* register *) pwire FA_cout_1797;
  (* register *) pwire FA_cout_1798;
  (* register *) pwire FA_cout_1799;
  (* register *) pwire FA_cout_1800;
  (* register *) pwire FA_cout_1801;
  (* register *) pwire FA_cout_1802;
  (* register *) pwire FA_cout_1803;
  (* register *) pwire FA_cout_1804;
  (* register *) pwire FA_cout_1805;
  (* register *) pwire FA_cout_1806;
  (* register *) pwire FA_cout_1807;
  (* register *) pwire FA_cout_1808;
  (* register *) pwire FA_cout_1809;
  (* register *) pwire FA_cout_1810;
  (* register *) pwire FA_cout_1811;
  (* register *) pwire FA_cout_1812;
  (* register *) pwire FA_cout_1813;
  (* register *) pwire FA_cout_1814;
  (* register *) pwire FA_cout_1815;
  (* register *) pwire FA_cout_1816;
  (* register *) pwire FA_cout_1817;
  (* register *) pwire FA_cout_1818;
  (* register *) pwire FA_cout_1819;
  (* register *) pwire FA_cout_1820;
  (* register *) pwire FA_cout_1821;
  (* register *) pwire FA_cout_1822;
  (* register *) pwire FA_cout_1823;
  (* register *) pwire FA_cout_1824;
  (* register *) pwire FA_cout_1825;
  (* register *) pwire FA_cout_1826;
  (* register *) pwire FA_cout_1827;
  (* register *) pwire FA_cout_1828;
  (* register *) pwire FA_cout_1829;
  (* register *) pwire FA_cout_1830;
  (* register *) pwire FA_cout_1831;
  (* register *) pwire FA_cout_1832;
  (* register *) pwire FA_cout_1833;
  (* register *) pwire FA_cout_1834;
  (* register *) pwire FA_cout_1835;
  (* register *) pwire FA_cout_1836;
  (* register *) pwire FA_cout_1837;
  (* register *) pwire FA_cout_1838;
  (* register *) pwire FA_cout_1839;
  (* register *) pwire FA_cout_1840;
  (* register *) pwire FA_cout_1841;
  (* register *) pwire FA_cout_1842;
  (* register *) pwire FA_cout_1843;
  (* register *) pwire FA_cout_1844;
  (* register *) pwire FA_cout_1845;
  (* register *) pwire FA_cout_1846;
  (* register *) pwire FA_cout_1847;
  (* register *) pwire FA_cout_1848;
  (* register *) pwire FA_cout_1849;
  (* register *) pwire FA_cout_1850;
  (* register *) pwire FA_cout_1851;
  (* register *) pwire FA_cout_1852;
  (* register *) pwire FA_cout_1853;
  (* register *) pwire FA_cout_1854;
  (* register *) pwire FA_cout_1855;
  (* register *) pwire FA_cout_1856;
  (* register *) pwire FA_cout_1857;
  (* register *) pwire FA_cout_1858;
  (* register *) pwire FA_cout_1859;
  (* register *) pwire FA_cout_1860;
  (* register *) pwire FA_cout_1861;
  (* register *) pwire FA_cout_1862;
  (* register *) pwire FA_cout_1863;
  (* register *) pwire FA_cout_1864;
  (* register *) pwire FA_cout_1865;
  (* register *) pwire FA_cout_1866;
  (* register *) pwire FA_cout_1867;
  (* register *) pwire FA_cout_1868;
  (* register *) pwire FA_cout_1869;
  (* register *) pwire FA_cout_1870;
  (* register *) pwire FA_cout_1871;
  (* register *) pwire FA_cout_1872;
  (* register *) pwire FA_cout_1873;
  (* register *) pwire FA_cout_1874;
  (* register *) pwire FA_cout_1875;
  (* register *) pwire FA_cout_1876;
  (* register *) pwire FA_cout_1877;
  (* register *) pwire FA_cout_1878;
  (* register *) pwire FA_cout_1879;
  (* register *) pwire FA_cout_1880;
  (* register *) pwire FA_cout_1881;
  (* register *) pwire FA_cout_1882;
  (* register *) pwire FA_cout_1883;
  (* register *) pwire FA_cout_1884;
  (* register *) pwire FA_cout_1885;
  (* register *) pwire FA_cout_1886;
  (* register *) pwire FA_cout_1887;
  (* register *) pwire FA_cout_1888;
  (* register *) pwire FA_cout_1889;
  (* register *) pwire FA_cout_1890;
  (* register *) pwire FA_cout_1891;
  (* register *) pwire FA_cout_1892;
  (* register *) pwire FA_cout_1893;
  (* register *) pwire FA_cout_1894;
  (* register *) pwire FA_cout_1895;
  (* register *) pwire FA_cout_1896;
  (* register *) pwire FA_cout_1897;
  (* register *) pwire FA_cout_1898;
  (* register *) pwire FA_cout_1899;
  (* register *) pwire FA_cout_1900;
  (* register *) pwire FA_cout_1901;
  (* register *) pwire FA_cout_1902;
  (* register *) pwire FA_cout_1903;
  (* register *) pwire FA_cout_1904;
  (* register *) pwire FA_cout_1905;
  (* register *) pwire FA_cout_1906;
  (* register *) pwire FA_cout_1907;
  (* register *) pwire FA_cout_1908;
  (* register *) pwire FA_cout_1909;
  (* register *) pwire FA_cout_1910;
  (* register *) pwire FA_cout_1911;
  (* register *) pwire FA_cout_1912;
  (* register *) pwire FA_cout_1913;
  (* register *) pwire FA_cout_1914;
  (* register *) pwire FA_cout_1915;
  (* register *) pwire FA_cout_1916;
  (* register *) pwire FA_cout_1917;
  (* register *) pwire FA_cout_1918;
  (* register *) pwire FA_cout_1919;
  (* register *) pwire FA_cout_1920;
  (* register *) pwire FA_cout_1921;
  (* register *) pwire FA_cout_1922;
  (* register *) pwire FA_cout_1923;
  (* register *) pwire FA_cout_1924;
  (* register *) pwire FA_cout_1925;
  (* register *) pwire FA_cout_1926;
  (* register *) pwire FA_cout_1927;
  (* register *) pwire FA_cout_1928;
  (* register *) pwire FA_cout_1929;
  (* register *) pwire FA_cout_1930;
  (* register *) pwire FA_cout_1931;
  (* register *) pwire FA_cout_1932;
  (* register *) pwire FA_cout_1933;
  (* register *) pwire FA_cout_1934;
  (* register *) pwire FA_cout_1935;
  (* register *) pwire FA_cout_1936;
  (* register *) pwire FA_cout_1937;
  (* register *) pwire FA_cout_1938;
  (* register *) pwire FA_cout_1939;
  (* register *) pwire FA_cout_1940;
  (* register *) pwire FA_cout_1941;
  (* register *) pwire FA_cout_1942;
  (* register *) pwire FA_cout_1943;
  (* register *) pwire FA_cout_1944;
  (* register *) pwire FA_cout_1945;
  (* register *) pwire FA_cout_1946;
  (* register *) pwire FA_cout_1947;
  (* register *) pwire FA_cout_1948;
  (* register *) pwire FA_cout_1949;
  (* register *) pwire FA_cout_1950;
  (* register *) pwire FA_cout_1951;
  (* register *) pwire FA_cout_1952;
  (* register *) pwire FA_cout_1953;
  (* register *) pwire FA_cout_1954;
  (* register *) pwire FA_cout_1955;
  (* register *) pwire FA_cout_1956;
  (* register *) pwire FA_cout_1957;
  (* register *) pwire FA_cout_1958;
  (* register *) pwire FA_cout_1959;
  (* register *) pwire FA_cout_1960;
  (* register *) pwire FA_cout_1961;
  (* register *) pwire FA_cout_1962;
  (* register *) pwire FA_cout_1963;
  (* register *) pwire FA_cout_1964;
  (* register *) pwire FA_cout_1965;
  (* register *) pwire FA_cout_1966;
  (* register *) pwire FA_cout_1967;
  (* register *) pwire FA_cout_1968;
  (* register *) pwire FA_cout_1969;
  (* register *) pwire FA_cout_1970;
  (* register *) pwire FA_cout_1971;
  (* register *) pwire FA_cout_1972;
  (* register *) pwire FA_cout_1973;
  (* register *) pwire FA_cout_1974;
  (* register *) pwire FA_cout_1975;
  (* register *) pwire FA_cout_1976;
  (* register *) pwire FA_cout_1977;
  (* register *) pwire FA_cout_1978;
  (* register *) pwire FA_cout_1979;
  (* register *) pwire FA_cout_1980;
  (* register *) pwire FA_cout_1981;
  (* register *) pwire FA_cout_1982;
  (* register *) pwire FA_cout_1983;
  (* register *) pwire FA_cout_1984;
  (* register *) pwire FA_cout_1985;
  (* register *) pwire FA_cout_1986;
  (* register *) pwire FA_cout_1987;
  (* register *) pwire FA_cout_1988;
  (* register *) pwire FA_cout_1989;
  (* register *) pwire FA_cout_1990;
  (* register *) pwire FA_cout_1991;
  (* register *) pwire FA_cout_1992;
  (* register *) pwire FA_cout_1993;
  (* register *) pwire FA_cout_1994;
  (* register *) pwire FA_cout_1995;
  (* register *) pwire FA_cout_1996;
  (* register *) pwire FA_cout_1997;
  (* register *) pwire FA_cout_1998;
  (* register *) pwire FA_cout_1999;
  (* register *) pwire FA_cout_2000;
  (* register *) pwire FA_cout_2001;
  (* register *) pwire FA_cout_2002;
  (* register *) pwire FA_cout_2003;
  (* register *) pwire FA_cout_2004;
  (* register *) pwire FA_cout_2005;
  (* register *) pwire FA_cout_2006;
  (* register *) pwire FA_cout_2007;
  (* register *) pwire FA_cout_2008;
  (* register *) pwire FA_cout_2009;
  (* register *) pwire FA_cout_2010;
  (* register *) pwire FA_cout_2011;
  (* register *) pwire FA_cout_2012;
  (* register *) pwire FA_cout_2013;
  (* register *) pwire FA_cout_2014;
  (* register *) pwire FA_cout_2015;
  (* register *) pwire FA_cout_2016;
  (* register *) pwire FA_cout_2017;
  (* register *) pwire FA_cout_2018;
  (* register *) pwire FA_cout_2019;
  (* register *) pwire FA_cout_2020;
  (* register *) pwire FA_cout_2021;
  (* register *) pwire FA_cout_2022;
  (* register *) pwire FA_cout_2023;
  (* register *) pwire FA_cout_2024;
  (* register *) pwire FA_cout_2025;
  (* register *) pwire FA_cout_2026;
  (* register *) pwire FA_cout_2027;
  (* register *) pwire FA_cout_2028;
  (* register *) pwire FA_cout_2029;
  (* register *) pwire FA_cout_2030;
  (* register *) pwire FA_cout_2031;
  (* register *) pwire FA_cout_2032;
  (* register *) pwire FA_cout_2033;
  (* register *) pwire FA_cout_2034;
  (* register *) pwire FA_cout_2035;
  (* register *) pwire FA_cout_2036;
  (* register *) pwire FA_cout_2037;
  (* register *) pwire FA_cout_2038;
  (* register *) pwire FA_cout_2039;
  (* register *) pwire FA_cout_2040;
  (* register *) pwire FA_cout_2041;
  (* register *) pwire FA_cout_2042;
  (* register *) pwire FA_cout_2043;
  (* register *) pwire FA_cout_2044;
  (* register *) pwire FA_cout_2045;
  (* register *) pwire FA_cout_2046;
  (* register *) pwire FA_cout_2047;
  (* register *) pwire FA_cout_2048;
  (* register *) pwire FA_cout_2049;
  (* register *) pwire FA_cout_2050;
  (* register *) pwire FA_cout_2051;
  (* register *) pwire FA_cout_2052;
  (* register *) pwire FA_cout_2053;
  (* register *) pwire FA_cout_2054;
  (* register *) pwire FA_cout_2055;
  (* register *) pwire FA_cout_2056;
  (* register *) pwire FA_cout_2057;
  (* register *) pwire FA_cout_2058;
  (* register *) pwire FA_cout_2059;
  (* register *) pwire FA_cout_2060;
  (* register *) pwire FA_cout_2061;
  (* register *) pwire FA_cout_2062;
  (* register *) pwire FA_cout_2063;
  (* register *) pwire FA_cout_2064;
  (* register *) pwire FA_cout_2065;
  (* register *) pwire FA_cout_2066;
  (* register *) pwire FA_cout_2067;
  (* register *) pwire FA_cout_2068;
  (* register *) pwire FA_cout_2069;
  (* register *) pwire FA_cout_2070;
  (* register *) pwire FA_cout_2071;
  (* register *) pwire FA_cout_2072;
  (* register *) pwire FA_cout_2073;
  (* register *) pwire FA_cout_2074;
  (* register *) pwire FA_cout_2075;
  (* register *) pwire FA_cout_2076;
  (* register *) pwire FA_cout_2077;
  (* register *) pwire FA_cout_2078;
  (* register *) pwire FA_cout_2079;
  (* register *) pwire FA_cout_2080;
  (* register *) pwire FA_cout_2081;
  (* register *) pwire FA_cout_2082;
  (* register *) pwire FA_cout_2083;
  (* register *) pwire FA_cout_2084;
  (* register *) pwire FA_cout_2085;
  (* register *) pwire FA_cout_2086;
  (* register *) pwire FA_cout_2087;
  (* register *) pwire FA_cout_2088;
  (* register *) pwire FA_cout_2089;
  (* register *) pwire FA_cout_2090;
  (* register *) pwire FA_cout_2091;
  (* register *) pwire FA_cout_2092;
  (* register *) pwire FA_cout_2093;
  (* register *) pwire FA_cout_2094;
  (* register *) pwire FA_cout_2095;
  (* register *) pwire FA_cout_2096;
  (* register *) pwire FA_cout_2097;
  (* register *) pwire FA_cout_2098;
  (* register *) pwire FA_cout_2099;
  (* register *) pwire FA_cout_2100;
  (* register *) pwire FA_cout_2101;
  (* register *) pwire FA_cout_2102;
  (* register *) pwire FA_cout_2103;
  (* register *) pwire FA_cout_2104;
  (* register *) pwire FA_cout_2105;
  (* register *) pwire FA_cout_2106;
  (* register *) pwire FA_cout_2107;
  (* register *) pwire FA_cout_2108;
  (* register *) pwire FA_cout_2109;
  (* register *) pwire FA_cout_2110;
  (* register *) pwire FA_cout_2111;
  (* register *) pwire FA_cout_2112;
  (* register *) pwire FA_cout_2113;
  (* register *) pwire FA_cout_2114;
  (* register *) pwire FA_cout_2115;
  (* register *) pwire FA_cout_2116;
  (* register *) pwire FA_cout_2117;
  (* register *) pwire FA_cout_2118;
  (* register *) pwire FA_cout_2119;
  (* register *) pwire FA_cout_2120;
  (* register *) pwire FA_cout_2121;
  (* register *) pwire FA_cout_2122;
  (* register *) pwire FA_cout_2123;
  (* register *) pwire FA_cout_2124;
  (* register *) pwire FA_cout_2125;
  (* register *) pwire FA_cout_2126;
  (* register *) pwire FA_cout_2127;
  (* register *) pwire FA_cout_2128;
  (* register *) pwire FA_cout_2129;
  (* register *) pwire FA_cout_2130;
  (* register *) pwire FA_cout_2131;
  (* register *) pwire FA_cout_2132;
  (* register *) pwire FA_cout_2133;
  (* register *) pwire FA_cout_2134;
  (* register *) pwire FA_cout_2135;
  (* register *) pwire FA_cout_2136;
  (* register *) pwire FA_cout_2137;
  (* register *) pwire FA_cout_2138;
  (* register *) pwire FA_cout_2139;
  (* register *) pwire FA_cout_2140;
  (* register *) pwire FA_cout_2141;
  (* register *) pwire FA_cout_2142;
  (* register *) pwire FA_cout_2143;
  (* register *) pwire FA_cout_2144;
  (* register *) pwire FA_cout_2145;
  (* register *) pwire FA_cout_2146;
  (* register *) pwire FA_cout_2147;
  (* register *) pwire FA_cout_2148;
  (* register *) pwire FA_cout_2149;
  (* register *) pwire FA_cout_2150;
  (* register *) pwire FA_cout_2151;
  (* register *) pwire FA_cout_2152;
  (* register *) pwire FA_cout_2153;
  (* register *) pwire FA_cout_2154;
  (* register *) pwire FA_cout_2155;
  (* register *) pwire FA_cout_2156;
  (* register *) pwire FA_cout_2157;
  (* register *) pwire FA_cout_2158;
  (* register *) pwire FA_cout_2159;
  (* register *) pwire FA_cout_2160;
  (* register *) pwire FA_cout_2161;
  (* register *) pwire FA_cout_2162;
  (* register *) pwire FA_cout_2163;
  (* register *) pwire FA_cout_2164;
  (* register *) pwire FA_cout_2165;
  (* register *) pwire FA_cout_2166;
  (* register *) pwire FA_cout_2167;
  (* register *) pwire FA_cout_2168;
  (* register *) pwire FA_cout_2169;
  (* register *) pwire FA_cout_2170;
  (* register *) pwire FA_cout_2171;
  (* register *) pwire FA_cout_2172;
  (* register *) pwire FA_cout_2173;
  (* register *) pwire FA_cout_2174;
  (* register *) pwire FA_cout_2175;
  (* register *) pwire FA_cout_2176;
  (* register *) pwire FA_cout_2177;
  (* register *) pwire FA_cout_2178;
  (* register *) pwire FA_cout_2179;
  (* register *) pwire FA_cout_2180;
  (* register *) pwire FA_cout_2181;
  (* register *) pwire FA_cout_2182;
  (* register *) pwire FA_cout_2183;
  (* register *) pwire FA_cout_2184;
  (* register *) pwire FA_cout_2185;
  (* register *) pwire FA_cout_2186;
  (* register *) pwire FA_cout_2187;
  (* register *) pwire FA_cout_2188;
  (* register *) pwire FA_cout_2189;
  (* register *) pwire FA_cout_2190;
  (* register *) pwire FA_cout_2191;
  (* register *) pwire FA_cout_2192;
  (* register *) pwire FA_cout_2193;
  (* register *) pwire FA_cout_2194;
  (* register *) pwire FA_cout_2195;
  (* register *) pwire FA_cout_2196;
  (* register *) pwire FA_cout_2197;
  (* register *) pwire FA_cout_2198;
  (* register *) pwire FA_cout_2199;
  (* register *) pwire FA_cout_2200;
  (* register *) pwire FA_cout_2201;
  (* register *) pwire FA_cout_2202;
  (* register *) pwire FA_cout_2203;
  (* register *) pwire FA_cout_2204;
  (* register *) pwire FA_cout_2205;
  (* register *) pwire FA_cout_2206;
  (* register *) pwire FA_cout_2207;
  (* register *) pwire FA_cout_2208;
  (* register *) pwire FA_cout_2209;
  (* register *) pwire FA_cout_2210;
  (* register *) pwire FA_cout_2211;
  (* register *) pwire FA_cout_2212;
  (* register *) pwire FA_cout_2213;
  (* register *) pwire FA_cout_2214;
  (* register *) pwire FA_cout_2215;
  (* register *) pwire FA_cout_2216;
  (* register *) pwire FA_cout_2217;
  (* register *) pwire FA_cout_2218;
  (* register *) pwire FA_cout_2219;
  (* register *) pwire FA_cout_2220;
  (* register *) pwire FA_cout_2221;
  (* register *) pwire FA_cout_2222;
  (* register *) pwire FA_cout_2223;
  (* register *) pwire FA_cout_2224;
  (* register *) pwire FA_cout_2225;
  (* register *) pwire FA_cout_2226;
  (* register *) pwire FA_cout_2227;
  (* register *) pwire FA_cout_2228;
  (* register *) pwire FA_cout_2229;
  (* register *) pwire FA_cout_2230;
  (* register *) pwire FA_cout_2231;
  (* register *) pwire FA_cout_2232;
  (* register *) pwire FA_cout_2233;
  (* register *) pwire FA_cout_2234;
  (* register *) pwire FA_cout_2235;
  (* register *) pwire FA_cout_2236;
  (* register *) pwire FA_cout_2237;
  (* register *) pwire FA_cout_2238;
  (* register *) pwire FA_cout_2239;
  (* register *) pwire FA_cout_2240;
  (* register *) pwire FA_cout_2241;
  (* register *) pwire FA_cout_2242;
  (* register *) pwire FA_cout_2243;
  (* register *) pwire FA_cout_2244;
  (* register *) pwire FA_cout_2245;
  (* register *) pwire FA_cout_2246;
  (* register *) pwire FA_cout_2247;
  (* register *) pwire FA_cout_2248;
  (* register *) pwire FA_cout_2249;
  (* register *) pwire FA_cout_2250;
  (* register *) pwire FA_cout_2251;
  (* register *) pwire FA_cout_2252;
  (* register *) pwire FA_cout_2253;
  (* register *) pwire FA_cout_2254;
  (* register *) pwire FA_cout_2255;
  (* register *) pwire FA_cout_2256;
  (* register *) pwire FA_cout_2257;
  (* register *) pwire FA_cout_2258;
  (* register *) pwire FA_cout_2259;
  (* register *) pwire FA_cout_2260;
  (* register *) pwire FA_cout_2261;
  (* register *) pwire FA_cout_2262;
  (* register *) pwire FA_cout_2263;
  (* register *) pwire FA_cout_2264;
  (* register *) pwire FA_cout_2265;
  (* register *) pwire FA_cout_2266;
  (* register *) pwire FA_cout_2267;
  (* register *) pwire FA_cout_2268;
  (* register *) pwire FA_cout_2269;
  (* register *) pwire FA_cout_2270;
  (* register *) pwire FA_cout_2271;
  (* register *) pwire FA_cout_2272;
  (* register *) pwire FA_cout_2273;
  (* register *) pwire FA_cout_2274;
  (* register *) pwire FA_cout_2275;
  (* register *) pwire FA_cout_2276;
  (* register *) pwire FA_cout_2277;
  (* register *) pwire FA_cout_2278;
  (* register *) pwire FA_cout_2279;
  (* register *) pwire FA_cout_2280;
  (* register *) pwire FA_cout_2281;
  (* register *) pwire FA_cout_2282;
  (* register *) pwire FA_cout_2283;
  (* register *) pwire FA_cout_2284;
  (* register *) pwire FA_cout_2285;
  (* register *) pwire FA_cout_2286;
  (* register *) pwire FA_cout_2287;
  (* register *) pwire FA_cout_2288;
  (* register *) pwire FA_cout_2289;
  (* register *) pwire FA_cout_2290;
  (* register *) pwire FA_cout_2291;
  (* register *) pwire FA_cout_2292;
  (* register *) pwire FA_cout_2293;
  (* register *) pwire FA_cout_2294;
  (* register *) pwire FA_cout_2295;
  (* register *) pwire FA_cout_2296;
  (* register *) pwire FA_cout_2297;
  (* register *) pwire FA_cout_2298;
  (* register *) pwire FA_cout_2299;
  (* register *) pwire FA_cout_2300;
  (* register *) pwire FA_cout_2301;
  (* register *) pwire FA_cout_2302;
  (* register *) pwire FA_cout_2303;
  (* register *) pwire FA_cout_2304;
  (* register *) pwire FA_cout_2305;
  (* register *) pwire FA_cout_2306;
  (* register *) pwire FA_cout_2307;
  (* register *) pwire FA_cout_2308;
  (* register *) pwire FA_cout_2309;
  (* register *) pwire FA_cout_2310;
  (* register *) pwire FA_cout_2311;
  (* register *) pwire FA_cout_2312;
  (* register *) pwire FA_cout_2313;
  (* register *) pwire FA_cout_2314;
  (* register *) pwire FA_cout_2315;
  (* register *) pwire FA_cout_2316;
  (* register *) pwire FA_cout_2317;
  (* register *) pwire FA_cout_2318;
  (* register *) pwire FA_cout_2319;
  (* register *) pwire FA_cout_2320;
  (* register *) pwire FA_cout_2321;
  (* register *) pwire FA_cout_2322;
  (* register *) pwire FA_cout_2323;
  (* register *) pwire FA_cout_2324;
  (* register *) pwire FA_cout_2325;
  (* register *) pwire FA_cout_2326;
  (* register *) pwire FA_cout_2327;
  (* register *) pwire FA_cout_2328;
  (* register *) pwire FA_cout_2329;
  (* register *) pwire FA_cout_2330;
  (* register *) pwire FA_cout_2331;
  (* register *) pwire FA_cout_2332;
  (* register *) pwire FA_cout_2333;
  (* register *) pwire FA_cout_2334;
  (* register *) pwire FA_cout_2335;
  (* register *) pwire FA_cout_2336;
  (* register *) pwire FA_cout_2337;
  (* register *) pwire FA_cout_2338;
  (* register *) pwire FA_cout_2339;
  (* register *) pwire FA_cout_2340;
  (* register *) pwire FA_cout_2341;
  (* register *) pwire FA_cout_2342;
  (* register *) pwire FA_cout_2343;
  (* register *) pwire FA_cout_2344;
  (* register *) pwire FA_cout_2345;
  (* register *) pwire FA_cout_2346;
  (* register *) pwire FA_cout_2347;
  (* register *) pwire FA_cout_2348;
  (* register *) pwire FA_cout_2349;
  (* register *) pwire FA_cout_2350;
  (* register *) pwire FA_cout_2351;
  (* register *) pwire FA_cout_2352;
  (* register *) pwire FA_cout_2353;
  (* register *) pwire FA_cout_2354;
  (* register *) pwire FA_cout_2355;
  (* register *) pwire FA_cout_2356;
  (* register *) pwire FA_cout_2357;
  (* register *) pwire FA_cout_2358;
  (* register *) pwire FA_cout_2359;
  (* register *) pwire FA_cout_2360;
  (* register *) pwire FA_cout_2361;
  (* register *) pwire FA_cout_2362;
  (* register *) pwire FA_cout_2363;
  (* register *) pwire FA_cout_2364;
  (* register *) pwire FA_cout_2365;
  (* register *) pwire FA_cout_2366;
  (* register *) pwire FA_cout_2367;
  (* register *) pwire FA_cout_2368;
  (* register *) pwire FA_cout_2369;
  (* register *) pwire FA_cout_2370;
  (* register *) pwire FA_cout_2371;
  (* register *) pwire FA_cout_2372;
  (* register *) pwire FA_cout_2373;
  (* register *) pwire FA_cout_2374;
  (* register *) pwire FA_cout_2375;
  (* register *) pwire FA_cout_2376;
  (* register *) pwire FA_cout_2377;
  (* register *) pwire FA_cout_2378;
  (* register *) pwire FA_cout_2379;
  (* register *) pwire FA_cout_2380;
  (* register *) pwire FA_cout_2381;
  (* register *) pwire FA_cout_2382;
  (* register *) pwire FA_cout_2383;
  (* register *) pwire FA_cout_2384;
  (* register *) pwire FA_cout_2385;
  (* register *) pwire FA_cout_2386;
  (* register *) pwire FA_cout_2387;
  (* register *) pwire FA_cout_2388;
  (* register *) pwire FA_cout_2389;
  (* register *) pwire FA_cout_2390;
  (* register *) pwire FA_cout_2391;
  (* register *) pwire FA_cout_2392;
  (* register *) pwire FA_cout_2393;
  (* register *) pwire FA_cout_2394;
  (* register *) pwire FA_cout_2395;
  (* register *) pwire FA_cout_2396;
  (* register *) pwire FA_cout_2397;
  (* register *) pwire FA_cout_2398;
  (* register *) pwire FA_cout_2399;
  (* register *) pwire FA_cout_2400;
  (* register *) pwire FA_cout_2401;
  (* register *) pwire FA_cout_2402;
  (* register *) pwire FA_cout_2403;
  (* register *) pwire FA_cout_2404;
  (* register *) pwire FA_cout_2405;
  (* register *) pwire FA_cout_2406;
  (* register *) pwire FA_cout_2407;
  (* register *) pwire FA_cout_2408;
  (* register *) pwire FA_cout_2409;
  (* register *) pwire FA_cout_2410;
  (* register *) pwire FA_cout_2411;
  (* register *) pwire FA_cout_2412;
  (* register *) pwire FA_cout_2413;
  (* register *) pwire FA_cout_2414;
  (* register *) pwire FA_cout_2415;
  (* register *) pwire FA_cout_2416;
  (* register *) pwire FA_cout_2417;
  (* register *) pwire FA_cout_2418;
  (* register *) pwire FA_cout_2419;
  (* register *) pwire FA_cout_2420;
  (* register *) pwire FA_cout_2421;
  (* register *) pwire FA_cout_2422;
  (* register *) pwire FA_cout_2423;
  (* register *) pwire FA_cout_2424;
  (* register *) pwire FA_cout_2425;
  (* register *) pwire FA_cout_2426;
  (* register *) pwire FA_cout_2427;
  (* register *) pwire FA_cout_2428;
  (* register *) pwire FA_cout_2429;
  (* register *) pwire FA_cout_2430;
  (* register *) pwire FA_cout_2431;
  (* register *) pwire FA_cout_2432;
  (* register *) pwire FA_cout_2433;
  (* register *) pwire FA_cout_2434;
  (* register *) pwire FA_cout_2435;
  (* register *) pwire FA_cout_2436;
  (* register *) pwire FA_cout_2437;
  (* register *) pwire FA_cout_2438;
  (* register *) pwire FA_cout_2439;
  (* register *) pwire FA_cout_2440;
  (* register *) pwire FA_cout_2441;
  (* register *) pwire FA_cout_2442;
  (* register *) pwire FA_cout_2443;
  (* register *) pwire FA_cout_2444;
  (* register *) pwire FA_cout_2445;
  (* register *) pwire FA_cout_2446;
  (* register *) pwire FA_cout_2447;
  (* register *) pwire FA_cout_2448;
  (* register *) pwire FA_cout_2449;
  (* register *) pwire FA_cout_2450;
  (* register *) pwire FA_cout_2451;
  (* register *) pwire FA_cout_2452;
  (* register *) pwire FA_cout_2453;
  (* register *) pwire FA_cout_2454;
  (* register *) pwire FA_cout_2455;
  (* register *) pwire FA_cout_2456;
  (* register *) pwire FA_cout_2457;
  (* register *) pwire FA_cout_2458;
  (* register *) pwire FA_cout_2459;
  (* register *) pwire FA_cout_2460;
  (* register *) pwire FA_cout_2461;
  (* register *) pwire FA_cout_2462;
  (* register *) pwire FA_cout_2463;
  (* register *) pwire FA_cout_2464;
  (* register *) pwire FA_cout_2465;
  (* register *) pwire FA_cout_2466;
  (* register *) pwire FA_cout_2467;
  (* register *) pwire FA_cout_2468;
  (* register *) pwire FA_cout_2469;
  (* register *) pwire FA_cout_2470;
  (* register *) pwire FA_cout_2471;
  (* register *) pwire FA_cout_2472;
  (* register *) pwire FA_cout_2473;
  (* register *) pwire FA_cout_2474;
  (* register *) pwire FA_cout_2475;
  (* register *) pwire FA_cout_2476;
  (* register *) pwire FA_cout_2477;
  (* register *) pwire FA_cout_2478;
  (* register *) pwire FA_cout_2479;
  (* register *) pwire FA_cout_2480;
  (* register *) pwire FA_cout_2481;
  (* register *) pwire FA_cout_2482;
  (* register *) pwire FA_cout_2483;
  (* register *) pwire FA_cout_2484;
  (* register *) pwire FA_cout_2485;
  (* register *) pwire FA_cout_2486;
  (* register *) pwire FA_cout_2487;
  (* register *) pwire FA_cout_2488;
  (* register *) pwire FA_cout_2489;
  (* register *) pwire FA_cout_2490;
  (* register *) pwire FA_cout_2491;
  (* register *) pwire FA_cout_2492;
  (* register *) pwire FA_cout_2493;
  (* register *) pwire FA_cout_2494;
  (* register *) pwire FA_cout_2495;
  (* register *) pwire FA_cout_2496;
  (* register *) pwire FA_cout_2497;
  (* register *) pwire FA_cout_2498;
  (* register *) pwire FA_cout_2499;
  (* register *) pwire FA_cout_2500;
  (* register *) pwire FA_cout_2501;
  (* register *) pwire FA_cout_2502;
  (* register *) pwire FA_cout_2503;
  (* register *) pwire FA_cout_2504;
  (* register *) pwire FA_cout_2505;
  (* register *) pwire FA_cout_2506;
  (* register *) pwire FA_cout_2507;
  (* register *) pwire FA_cout_2508;
  (* register *) pwire FA_cout_2509;
  (* register *) pwire FA_cout_2510;
  (* register *) pwire FA_cout_2511;
  (* register *) pwire FA_cout_2512;
  (* register *) pwire FA_cout_2513;
  (* register *) pwire FA_cout_2514;
  (* register *) pwire FA_cout_2515;
  (* register *) pwire FA_cout_2516;
  (* register *) pwire FA_cout_2517;
  (* register *) pwire FA_cout_2518;
  (* register *) pwire FA_cout_2519;
  (* register *) pwire FA_cout_2520;
  (* register *) pwire FA_cout_2521;
  (* register *) pwire FA_cout_2522;
  (* register *) pwire FA_cout_2523;
  (* register *) pwire FA_cout_2524;
  (* register *) pwire FA_cout_2525;
  (* register *) pwire FA_cout_2526;
  (* register *) pwire FA_cout_2527;
  (* register *) pwire FA_cout_2528;
  (* register *) pwire FA_cout_2529;
  (* register *) pwire FA_cout_2530;
  (* register *) pwire FA_cout_2531;
  (* register *) pwire FA_cout_2532;
  (* register *) pwire FA_cout_2533;
  (* register *) pwire FA_cout_2534;
  (* register *) pwire FA_cout_2535;
  (* register *) pwire FA_cout_2536;
  (* register *) pwire FA_cout_2537;
  (* register *) pwire FA_cout_2538;
  (* register *) pwire FA_cout_2539;
  (* register *) pwire FA_cout_2540;
  (* register *) pwire FA_cout_2541;
  (* register *) pwire FA_cout_2542;
  (* register *) pwire FA_cout_2543;
  (* register *) pwire FA_cout_2544;
  (* register *) pwire FA_cout_2545;
  (* register *) pwire FA_cout_2546;
  (* register *) pwire FA_cout_2547;
  (* register *) pwire FA_cout_2548;
  (* register *) pwire FA_cout_2549;
  (* register *) pwire FA_cout_2550;
  (* register *) pwire FA_cout_2551;
  (* register *) pwire FA_cout_2552;
  (* register *) pwire FA_cout_2553;
  (* register *) pwire FA_cout_2554;
  (* register *) pwire FA_cout_2555;
  (* register *) pwire FA_cout_2556;
  (* register *) pwire FA_cout_2557;
  (* register *) pwire FA_cout_2558;
  (* register *) pwire FA_cout_2559;
  (* register *) pwire FA_cout_2560;
  (* register *) pwire FA_cout_2561;
  (* register *) pwire FA_cout_2562;
  (* register *) pwire FA_cout_2563;
  (* register *) pwire FA_cout_2564;
  (* register *) pwire FA_cout_2565;
  (* register *) pwire FA_cout_2566;
  (* register *) pwire FA_cout_2567;
  (* register *) pwire FA_cout_2568;
  (* register *) pwire FA_cout_2569;
  (* register *) pwire FA_cout_2570;
  (* register *) pwire FA_cout_2571;
  (* register *) pwire FA_cout_2572;
  (* register *) pwire FA_cout_2573;
  (* register *) pwire FA_cout_2574;
  (* register *) pwire FA_cout_2575;
  (* register *) pwire FA_cout_2576;
  (* register *) pwire FA_cout_2577;
  (* register *) pwire FA_cout_2578;
  (* register *) pwire FA_cout_2579;
  (* register *) pwire FA_cout_2580;
  (* register *) pwire FA_cout_2581;
  (* register *) pwire FA_cout_2582;
  (* register *) pwire FA_cout_2583;
  (* register *) pwire FA_cout_2584;
  (* register *) pwire FA_cout_2585;
  (* register *) pwire FA_cout_2586;
  (* register *) pwire FA_cout_2587;
  (* register *) pwire FA_cout_2588;
  (* register *) pwire FA_cout_2589;
  (* register *) pwire FA_cout_2590;
  (* register *) pwire FA_cout_2591;
  (* register *) pwire FA_cout_2592;
  (* register *) pwire FA_cout_2593;
  (* register *) pwire FA_cout_2594;
  (* register *) pwire FA_cout_2595;
  (* register *) pwire FA_cout_2596;
  (* register *) pwire FA_cout_2597;
  (* register *) pwire FA_cout_2598;
  (* register *) pwire FA_cout_2599;
  (* register *) pwire FA_cout_2600;
  (* register *) pwire FA_cout_2601;
  (* register *) pwire FA_cout_2602;
  (* register *) pwire FA_cout_2603;
  (* register *) pwire FA_cout_2604;
  (* register *) pwire FA_cout_2605;
  (* register *) pwire FA_cout_2606;
  (* register *) pwire FA_cout_2607;
  (* register *) pwire FA_cout_2608;
  (* register *) pwire FA_cout_2609;
  (* register *) pwire FA_cout_2610;
  (* register *) pwire FA_cout_2611;
  (* register *) pwire FA_cout_2612;
  (* register *) pwire FA_cout_2613;
  (* register *) pwire FA_cout_2614;
  (* register *) pwire FA_cout_2615;
  (* register *) pwire FA_cout_2616;
  (* register *) pwire FA_cout_2617;
  (* register *) pwire FA_cout_2618;
  (* register *) pwire FA_cout_2619;
  (* register *) pwire FA_cout_2620;
  (* register *) pwire FA_cout_2621;
  (* register *) pwire FA_cout_2622;
  (* register *) pwire FA_cout_2623;
  (* register *) pwire FA_cout_2624;
  (* register *) pwire FA_cout_2625;
  (* register *) pwire FA_cout_2626;
  (* register *) pwire FA_cout_2627;
  (* register *) pwire FA_cout_2628;
  (* register *) pwire FA_cout_2629;
  (* register *) pwire FA_cout_2630;
  (* register *) pwire FA_cout_2631;
  (* register *) pwire FA_cout_2632;
  (* register *) pwire FA_cout_2633;
  (* register *) pwire FA_cout_2634;
  (* register *) pwire FA_cout_2635;
  (* register *) pwire FA_cout_2636;
  (* register *) pwire FA_cout_2637;
  (* register *) pwire FA_cout_2638;
  (* register *) pwire FA_cout_2639;
  (* register *) pwire FA_cout_2640;
  (* register *) pwire FA_cout_2641;
  (* register *) pwire FA_cout_2642;
  (* register *) pwire FA_cout_2643;
  (* register *) pwire FA_cout_2644;
  (* register *) pwire FA_cout_2645;
  (* register *) pwire FA_cout_2646;
  (* register *) pwire FA_cout_2647;
  (* register *) pwire FA_cout_2648;
  (* register *) pwire FA_cout_2649;
  (* register *) pwire FA_cout_2650;
  (* register *) pwire FA_cout_2651;
  (* register *) pwire FA_cout_2652;
  (* register *) pwire FA_cout_2653;
  (* register *) pwire FA_cout_2654;
  (* register *) pwire FA_cout_2655;
  (* register *) pwire FA_cout_2656;
  (* register *) pwire FA_cout_2657;
  (* register *) pwire FA_cout_2658;
  (* register *) pwire FA_cout_2659;
  (* register *) pwire FA_cout_2660;
  (* register *) pwire FA_cout_2661;
  (* register *) pwire FA_cout_2662;
  (* register *) pwire FA_cout_2663;
  (* register *) pwire FA_cout_2664;
  (* register *) pwire FA_cout_2665;
  (* register *) pwire FA_cout_2666;
  (* register *) pwire FA_cout_2667;
  (* register *) pwire FA_cout_2668;
  (* register *) pwire FA_cout_2669;
  (* register *) pwire FA_cout_2670;
  (* register *) pwire FA_cout_2671;
  (* register *) pwire FA_cout_2672;
  (* register *) pwire FA_cout_2673;
  (* register *) pwire FA_cout_2674;
  (* register *) pwire FA_cout_2675;
  (* register *) pwire FA_cout_2676;
  (* register *) pwire FA_cout_2677;
  (* register *) pwire FA_cout_2678;
  (* register *) pwire FA_cout_2679;
  (* register *) pwire FA_cout_2680;
  (* register *) pwire FA_cout_2681;
  (* register *) pwire FA_cout_2682;
  (* register *) pwire FA_cout_2683;
  (* register *) pwire FA_cout_2684;
  (* register *) pwire FA_cout_2685;
  (* register *) pwire FA_cout_2686;
  (* register *) pwire FA_cout_2687;
  (* register *) pwire FA_cout_2688;
  (* register *) pwire FA_cout_2689;
  (* register *) pwire FA_cout_2690;
  (* register *) pwire FA_cout_2691;
  (* register *) pwire FA_cout_2692;
  (* register *) pwire FA_cout_2693;
  (* register *) pwire FA_cout_2694;
  (* register *) pwire FA_cout_2695;
  (* register *) pwire FA_cout_2696;
  (* register *) pwire FA_cout_2697;
  (* register *) pwire FA_cout_2698;
  (* register *) pwire FA_cout_2699;
  (* register *) pwire FA_cout_2700;
  (* register *) pwire FA_cout_2701;
  (* register *) pwire FA_cout_2702;
  (* register *) pwire FA_cout_2703;
  (* register *) pwire FA_cout_2704;
  (* register *) pwire FA_cout_2705;
  (* register *) pwire FA_cout_2706;
  (* register *) pwire FA_cout_2707;
  (* register *) pwire FA_cout_2708;
  (* register *) pwire FA_cout_2709;
  (* register *) pwire FA_cout_2710;
  (* register *) pwire FA_cout_2711;
  (* register *) pwire FA_cout_2712;
  (* register *) pwire FA_cout_2713;
  (* register *) pwire FA_cout_2714;
  (* register *) pwire FA_cout_2715;
  (* register *) pwire FA_cout_2716;
  (* register *) pwire FA_cout_2717;
  (* register *) pwire FA_cout_2718;
  (* register *) pwire FA_cout_2719;
  (* register *) pwire FA_cout_2720;
  (* register *) pwire FA_cout_2721;
  (* register *) pwire FA_cout_2722;
  (* register *) pwire FA_cout_2723;
  (* register *) pwire FA_cout_2724;
  (* register *) pwire FA_cout_2725;
  (* register *) pwire FA_cout_2726;
  (* register *) pwire FA_cout_2727;
  (* register *) pwire FA_cout_2728;
  (* register *) pwire FA_cout_2729;
  (* register *) pwire FA_cout_2730;
  (* register *) pwire FA_cout_2731;
  (* register *) pwire FA_cout_2732;
  (* register *) pwire FA_cout_2733;
  (* register *) pwire FA_cout_2734;
  (* register *) pwire FA_cout_2735;
  (* register *) pwire FA_cout_2736;
  (* register *) pwire FA_cout_2737;
  (* register *) pwire FA_cout_2738;
  (* register *) pwire FA_cout_2739;
  (* register *) pwire FA_cout_2740;
  (* register *) pwire FA_cout_2741;
  (* register *) pwire FA_cout_2742;
  (* register *) pwire FA_cout_2743;
  (* register *) pwire FA_cout_2744;
  (* register *) pwire FA_cout_2745;
  (* register *) pwire FA_cout_2746;
  (* register *) pwire FA_cout_2747;
  (* register *) pwire FA_cout_2748;
  (* register *) pwire FA_cout_2749;
  (* register *) pwire FA_cout_2750;
  (* register *) pwire FA_cout_2751;
  (* register *) pwire FA_cout_2752;
  (* register *) pwire FA_cout_2753;
  (* register *) pwire FA_cout_2754;
  (* register *) pwire FA_cout_2755;
  (* register *) pwire FA_cout_2756;
  (* register *) pwire FA_cout_2757;
  (* register *) pwire FA_cout_2758;
  (* register *) pwire FA_cout_2759;
  (* register *) pwire FA_cout_2760;
  (* register *) pwire FA_cout_2761;
  (* register *) pwire FA_cout_2762;
  (* register *) pwire FA_cout_2763;
  (* register *) pwire FA_cout_2764;
  (* register *) pwire FA_cout_2765;
  (* register *) pwire FA_cout_2766;
  (* register *) pwire FA_cout_2767;
  (* register *) pwire FA_cout_2768;
  (* register *) pwire FA_cout_2769;
  (* register *) pwire FA_cout_2770;
  (* register *) pwire FA_cout_2771;
  (* register *) pwire FA_cout_2772;
  (* register *) pwire FA_cout_2773;
  (* register *) pwire FA_cout_2774;
  (* register *) pwire FA_cout_2775;
  (* register *) pwire FA_cout_2776;
  (* register *) pwire FA_cout_2777;
  (* register *) pwire FA_cout_2778;
  (* register *) pwire FA_cout_2779;
  (* register *) pwire FA_cout_2780;
  (* register *) pwire FA_cout_2781;
  (* register *) pwire FA_cout_2782;
  (* register *) pwire FA_cout_2783;
  (* register *) pwire FA_cout_2784;
  (* register *) pwire FA_cout_2785;
  (* register *) pwire FA_cout_2786;
  (* register *) pwire FA_cout_2787;
  (* register *) pwire FA_cout_2788;
  (* register *) pwire FA_cout_2789;
  (* register *) pwire FA_cout_2790;
  (* register *) pwire FA_cout_2791;
  (* register *) pwire FA_cout_2792;
  (* register *) pwire FA_cout_2793;
  (* register *) pwire FA_cout_2794;
  (* register *) pwire FA_cout_2795;
  (* register *) pwire FA_cout_2796;
  (* register *) pwire FA_cout_2797;
  (* register *) pwire FA_cout_2798;
  (* register *) pwire FA_cout_2799;
  (* register *) pwire FA_cout_2800;
  (* register *) pwire FA_cout_2801;
  (* register *) pwire FA_cout_2802;
  (* register *) pwire FA_cout_2803;
  (* register *) pwire FA_cout_2804;
  (* register *) pwire FA_cout_2805;
  (* register *) pwire FA_cout_2806;
  (* register *) pwire FA_cout_2807;
  (* register *) pwire FA_cout_2808;
  (* register *) pwire FA_cout_2809;
  (* register *) pwire FA_cout_2810;
  (* register *) pwire FA_cout_2811;
  (* register *) pwire FA_cout_2812;
  (* register *) pwire FA_cout_2813;
  (* register *) pwire FA_cout_2814;
  (* register *) pwire FA_cout_2815;
  (* register *) pwire FA_cout_2816;
  (* register *) pwire FA_cout_2817;
  (* register *) pwire FA_cout_2818;
  (* register *) pwire FA_cout_2819;
  (* register *) pwire FA_cout_2820;
  (* register *) pwire FA_cout_2821;
  (* register *) pwire FA_cout_2822;
  (* register *) pwire FA_cout_2823;
  (* register *) pwire FA_cout_2824;
  (* register *) pwire FA_cout_2825;
  (* register *) pwire FA_cout_2826;
  (* register *) pwire FA_cout_2827;
  (* register *) pwire FA_cout_2828;
  (* register *) pwire FA_cout_2829;
  (* register *) pwire FA_cout_2830;
  (* register *) pwire FA_cout_2831;
  (* register *) pwire FA_cout_2832;
  (* register *) pwire FA_cout_2833;
  (* register *) pwire FA_cout_2834;
  (* register *) pwire FA_cout_2835;
  (* register *) pwire FA_cout_2836;
  (* register *) pwire FA_cout_2837;
  (* register *) pwire FA_cout_2838;
  (* register *) pwire FA_cout_2839;
  (* register *) pwire FA_cout_2840;
  (* register *) pwire FA_cout_2841;
  (* register *) pwire FA_cout_2842;
  (* register *) pwire FA_cout_2843;
  (* register *) pwire FA_cout_2844;
  (* register *) pwire FA_cout_2845;
  (* register *) pwire FA_cout_2846;
  (* register *) pwire FA_cout_2847;
  (* register *) pwire FA_cout_2848;
  (* register *) pwire FA_cout_2849;
  (* register *) pwire FA_cout_2850;
  (* register *) pwire FA_cout_2851;
  (* register *) pwire FA_cout_2852;
  (* register *) pwire FA_cout_2853;
  (* register *) pwire FA_cout_2854;
  (* register *) pwire FA_cout_2855;
  (* register *) pwire FA_cout_2856;
  (* register *) pwire FA_cout_2857;
  (* register *) pwire FA_cout_2858;
  (* register *) pwire FA_cout_2859;
  (* register *) pwire FA_cout_2860;
  (* register *) pwire FA_cout_2861;
  (* register *) pwire FA_cout_2862;
  (* register *) pwire FA_cout_2863;
  (* register *) pwire FA_cout_2864;
  (* register *) pwire FA_cout_2865;
  (* register *) pwire FA_cout_2866;
  (* register *) pwire FA_cout_2867;
  (* register *) pwire FA_cout_2868;
  (* register *) pwire FA_cout_2869;
  (* register *) pwire FA_cout_2870;
  (* register *) pwire FA_cout_2871;
  (* register *) pwire FA_cout_2872;
  (* register *) pwire FA_cout_2873;
  (* register *) pwire FA_cout_2874;
  (* register *) pwire FA_cout_2875;
  (* register *) pwire FA_cout_2876;
  (* register *) pwire FA_cout_2877;
  (* register *) pwire FA_cout_2878;
  (* register *) pwire FA_cout_2879;
  (* register *) pwire FA_cout_2880;
  (* register *) pwire FA_cout_2881;
  (* register *) pwire FA_cout_2882;
  (* register *) pwire FA_cout_2883;
  (* register *) pwire FA_cout_2884;
  (* register *) pwire FA_cout_2885;
  (* register *) pwire FA_cout_2886;
  (* register *) pwire FA_cout_2887;
  (* register *) pwire FA_cout_2888;
  (* register *) pwire FA_cout_2889;
  (* register *) pwire FA_cout_2890;
  (* register *) pwire FA_cout_2891;
  (* register *) pwire FA_cout_2892;
  (* register *) pwire FA_cout_2893;
  (* register *) pwire FA_cout_2894;
  (* register *) pwire FA_cout_2895;
  (* register *) pwire FA_cout_2896;
  (* register *) pwire FA_cout_2897;
  (* register *) pwire FA_cout_2898;
  (* register *) pwire FA_cout_2899;
  (* register *) pwire FA_cout_2900;
  (* register *) pwire FA_cout_2901;
  (* register *) pwire FA_cout_2902;
  (* register *) pwire FA_cout_2903;
  (* register *) pwire FA_cout_2904;
  (* register *) pwire FA_cout_2905;
  (* register *) pwire FA_cout_2906;
  (* register *) pwire FA_cout_2907;
  (* register *) pwire FA_cout_2908;
  (* register *) pwire FA_cout_2909;
  (* register *) pwire FA_cout_2910;
  (* register *) pwire FA_cout_2911;
  (* register *) pwire FA_cout_2912;
  (* register *) pwire FA_cout_2913;
  (* register *) pwire FA_cout_2914;
  (* register *) pwire FA_cout_2915;
  (* register *) pwire FA_cout_2916;
  (* register *) pwire FA_cout_2917;
  (* register *) pwire FA_cout_2918;
  (* register *) pwire FA_cout_2919;
  (* register *) pwire FA_cout_2920;
  (* register *) pwire FA_cout_2921;
  (* register *) pwire FA_cout_2922;
  (* register *) pwire FA_cout_2923;
  (* register *) pwire FA_cout_2924;
  (* register *) pwire FA_cout_2925;
  (* register *) pwire FA_cout_2926;
  (* register *) pwire FA_cout_2927;
  (* register *) pwire FA_cout_2928;
  (* register *) pwire FA_cout_2929;
  (* register *) pwire FA_cout_2930;
  (* register *) pwire FA_cout_2931;
  (* register *) pwire FA_cout_2932;
  (* register *) pwire FA_cout_2933;
  (* register *) pwire FA_cout_2934;
  (* register *) pwire FA_cout_2935;
  (* register *) pwire FA_cout_2936;
  (* register *) pwire FA_cout_2937;
  (* register *) pwire FA_cout_2938;
  (* register *) pwire FA_cout_2939;
  (* register *) pwire FA_cout_2940;
  (* register *) pwire FA_cout_2941;
  (* register *) pwire FA_cout_2942;
  (* register *) pwire FA_cout_2943;
  (* register *) pwire FA_cout_2944;
  (* register *) pwire FA_cout_2945;
  (* register *) pwire FA_cout_2946;
  (* register *) pwire FA_cout_2947;
  (* register *) pwire FA_cout_2948;
  (* register *) pwire FA_cout_2949;
  (* register *) pwire FA_cout_2950;
  (* register *) pwire FA_cout_2951;
  (* register *) pwire FA_cout_2952;
  (* register *) pwire FA_cout_2953;
  (* register *) pwire FA_cout_2954;
  (* register *) pwire FA_cout_2955;
  (* register *) pwire FA_cout_2956;
  (* register *) pwire FA_cout_2957;
  (* register *) pwire FA_cout_2958;
  (* register *) pwire FA_cout_2959;
  (* register *) pwire FA_cout_2960;
  (* register *) pwire FA_cout_2961;
  (* register *) pwire FA_cout_2962;
  (* register *) pwire FA_cout_2963;
  (* register *) pwire FA_cout_2964;
  (* register *) pwire FA_cout_2965;
  (* register *) pwire FA_cout_2966;
  (* register *) pwire FA_cout_2967;
  (* register *) pwire FA_cout_2968;
  (* register *) pwire FA_cout_2969;
  (* register *) pwire FA_cout_2970;
  (* register *) pwire FA_cout_2971;
  (* register *) pwire FA_cout_2972;
  (* register *) pwire FA_cout_2973;
  (* register *) pwire FA_cout_2974;
  (* register *) pwire FA_cout_2975;
  (* register *) pwire FA_cout_2976;
  (* register *) pwire FA_cout_2977;
  (* register *) pwire FA_cout_2978;
  (* register *) pwire FA_cout_2979;
  (* register *) pwire FA_cout_2980;
  (* register *) pwire FA_cout_2981;
  (* register *) pwire FA_cout_2982;
  (* register *) pwire FA_cout_2983;
  (* register *) pwire FA_cout_2984;
  (* register *) pwire FA_cout_2985;
  (* register *) pwire FA_cout_2986;
  (* register *) pwire FA_cout_2987;
  (* register *) pwire FA_cout_2988;
  (* register *) pwire FA_cout_2989;
  (* register *) pwire FA_cout_2990;
  (* register *) pwire FA_cout_2991;
  (* register *) pwire FA_cout_2992;
  (* register *) pwire FA_cout_2993;
  (* register *) pwire FA_cout_2994;
  (* register *) pwire FA_cout_2995;
  (* register *) pwire FA_cout_2996;
  (* register *) pwire FA_cout_2997;
  (* register *) pwire FA_cout_2998;
  (* register *) pwire FA_cout_2999;
  (* register *) pwire FA_cout_3000;
  (* register *) pwire FA_cout_3001;
  (* register *) pwire FA_cout_3002;
  (* register *) pwire FA_cout_3003;
  (* register *) pwire FA_cout_3004;
  (* register *) pwire FA_cout_3005;
  (* register *) pwire FA_cout_3006;
  (* register *) pwire FA_cout_3007;
  (* register *) pwire FA_cout_3008;
  (* register *) pwire FA_cout_3009;
  (* register *) pwire FA_cout_3010;
  (* register *) pwire FA_cout_3011;
  (* register *) pwire FA_cout_3012;
  (* register *) pwire FA_cout_3013;
  (* register *) pwire FA_cout_3014;
  (* register *) pwire FA_cout_3015;
  (* register *) pwire FA_cout_3016;
  (* register *) pwire FA_cout_3017;
  (* register *) pwire FA_cout_3018;
  (* register *) pwire FA_cout_3019;
  (* register *) pwire FA_cout_3020;
  (* register *) pwire FA_cout_3021;
  (* register *) pwire FA_cout_3022;
  (* register *) pwire FA_cout_3023;
  (* register *) pwire FA_cout_3024;
  (* register *) pwire FA_cout_3025;
  (* register *) pwire FA_cout_3026;
  (* register *) pwire FA_cout_3027;
  (* register *) pwire FA_cout_3028;
  (* register *) pwire FA_cout_3029;
  (* register *) pwire FA_cout_3030;
  (* register *) pwire FA_cout_3031;
  (* register *) pwire FA_cout_3032;
  (* register *) pwire FA_cout_3033;
  (* register *) pwire FA_cout_3034;
  (* register *) pwire FA_cout_3035;
  (* register *) pwire FA_cout_3036;
  (* register *) pwire FA_cout_3037;
  (* register *) pwire FA_cout_3038;
  (* register *) pwire FA_cout_3039;
  (* register *) pwire FA_cout_3040;
  (* register *) pwire FA_cout_3041;
  (* register *) pwire FA_cout_3042;
  (* register *) pwire FA_cout_3043;
  (* register *) pwire FA_cout_3044;
  (* register *) pwire FA_cout_3045;
  (* register *) pwire FA_cout_3046;
  (* register *) pwire FA_cout_3047;
  (* register *) pwire FA_cout_3048;
  (* register *) pwire FA_cout_3049;
  (* register *) pwire FA_cout_3050;
  (* register *) pwire FA_cout_3051;
  (* register *) pwire FA_cout_3052;
  (* register *) pwire FA_cout_3053;
  (* register *) pwire FA_cout_3054;
  (* register *) pwire FA_cout_3055;
  (* register *) pwire FA_cout_3056;
  (* register *) pwire FA_cout_3057;
  (* register *) pwire FA_cout_3058;
  (* register *) pwire FA_cout_3059;
  (* register *) pwire FA_cout_3060;
  (* register *) pwire FA_cout_3061;
  (* register *) pwire FA_cout_3062;
  (* register *) pwire FA_cout_3063;
  (* register *) pwire FA_cout_3064;
  (* register *) pwire FA_cout_3065;
  (* register *) pwire FA_cout_3066;
  (* register *) pwire FA_cout_3067;
  (* register *) pwire FA_cout_3068;
  (* register *) pwire FA_cout_3069;
  (* register *) pwire FA_cout_3070;
  (* register *) pwire FA_cout_3071;
  (* register *) pwire FA_cout_3072;
  (* register *) pwire FA_cout_3073;
  (* register *) pwire FA_cout_3074;
  (* register *) pwire FA_cout_3075;
  (* register *) pwire FA_cout_3076;
  (* register *) pwire FA_cout_3077;
  (* register *) pwire FA_cout_3078;
  (* register *) pwire FA_cout_3079;
  (* register *) pwire FA_cout_3080;
  (* register *) pwire FA_cout_3081;
  (* register *) pwire FA_cout_3082;
  (* register *) pwire FA_cout_3083;
  (* register *) pwire FA_cout_3084;
  (* register *) pwire FA_cout_3085;
  (* register *) pwire FA_cout_3086;
  (* register *) pwire FA_cout_3087;
  (* register *) pwire FA_cout_3088;
  (* register *) pwire FA_cout_3089;
  (* register *) pwire FA_cout_3090;
  (* register *) pwire FA_cout_3091;
  (* register *) pwire FA_cout_3092;
  (* register *) pwire FA_cout_3093;
  (* register *) pwire FA_cout_3094;
  (* register *) pwire FA_cout_3095;
  (* register *) pwire FA_cout_3096;
  (* register *) pwire FA_cout_3097;
  (* register *) pwire FA_cout_3098;
  (* register *) pwire FA_cout_3099;
  (* register *) pwire FA_cout_3100;
  (* register *) pwire FA_cout_3101;
  (* register *) pwire FA_cout_3102;
  (* register *) pwire FA_cout_3103;
  (* register *) pwire FA_cout_3104;
  (* register *) pwire FA_cout_3105;
  (* register *) pwire FA_cout_3106;
  (* register *) pwire FA_cout_3107;
  (* register *) pwire FA_cout_3108;
  (* register *) pwire FA_cout_3109;
  (* register *) pwire FA_cout_3110;
  (* register *) pwire FA_cout_3111;
  (* register *) pwire FA_cout_3112;
  (* register *) pwire FA_cout_3113;
  (* register *) pwire FA_cout_3114;
  (* register *) pwire FA_cout_3115;
  (* register *) pwire FA_cout_3116;
  (* register *) pwire FA_cout_3117;
  (* register *) pwire FA_cout_3118;
  (* register *) pwire FA_cout_3119;
  (* register *) pwire FA_cout_3120;
  (* register *) pwire FA_cout_3121;
  (* register *) pwire FA_cout_3122;
  (* register *) pwire FA_cout_3123;
  (* register *) pwire FA_cout_3124;
  (* register *) pwire FA_cout_3125;
  (* register *) pwire FA_cout_3126;
  (* register *) pwire FA_cout_3127;
  (* register *) pwire FA_cout_3128;
  (* register *) pwire FA_cout_3129;
  (* register *) pwire FA_cout_3130;
  (* register *) pwire FA_cout_3131;
  (* register *) pwire FA_cout_3132;
  (* register *) pwire FA_cout_3133;
  (* register *) pwire FA_cout_3134;
  (* register *) pwire FA_cout_3135;
  (* register *) pwire FA_cout_3136;
  (* register *) pwire FA_cout_3137;
  (* register *) pwire FA_cout_3138;
  (* register *) pwire FA_cout_3139;
  (* register *) pwire FA_cout_3140;
  (* register *) pwire FA_cout_3141;
  (* register *) pwire FA_cout_3142;
  (* register *) pwire FA_cout_3143;
  (* register *) pwire FA_cout_3144;
  (* register *) pwire FA_cout_3145;
  (* register *) pwire FA_cout_3146;
  (* register *) pwire FA_cout_3147;
  (* register *) pwire FA_cout_3148;
  (* register *) pwire FA_cout_3149;
  (* register *) pwire FA_cout_3150;
  (* register *) pwire FA_cout_3151;
  (* register *) pwire FA_cout_3152;
  (* register *) pwire FA_cout_3153;
  (* register *) pwire FA_cout_3154;
  (* register *) pwire FA_cout_3155;
  (* register *) pwire FA_cout_3156;
  (* register *) pwire FA_cout_3157;
  (* register *) pwire FA_cout_3158;
  (* register *) pwire FA_cout_3159;
  (* register *) pwire FA_cout_3160;
  (* register *) pwire FA_cout_3161;
  (* register *) pwire FA_cout_3162;
  (* register *) pwire FA_cout_3163;
  (* register *) pwire FA_cout_3164;
  (* register *) pwire FA_cout_3165;
  (* register *) pwire FA_cout_3166;
  (* register *) pwire FA_cout_3167;
  (* register *) pwire FA_cout_3168;
  (* register *) pwire FA_cout_3169;
  (* register *) pwire FA_cout_3170;
  (* register *) pwire FA_cout_3171;
  (* register *) pwire FA_cout_3172;
  (* register *) pwire FA_cout_3173;
  (* register *) pwire FA_cout_3174;
  (* register *) pwire FA_cout_3175;
  (* register *) pwire FA_cout_3176;
  (* register *) pwire FA_cout_3177;
  (* register *) pwire FA_cout_3178;
  (* register *) pwire FA_cout_3179;
  (* register *) pwire FA_cout_3180;
  (* register *) pwire FA_cout_3181;
  (* register *) pwire FA_cout_3182;
  (* register *) pwire FA_cout_3183;
  (* register *) pwire FA_cout_3184;
  (* register *) pwire FA_cout_3185;
  (* register *) pwire FA_cout_3186;
  (* register *) pwire FA_cout_3187;
  (* register *) pwire FA_cout_3188;
  (* register *) pwire FA_cout_3189;
  (* register *) pwire FA_cout_3190;
  (* register *) pwire FA_cout_3191;
  (* register *) pwire FA_cout_3192;
  (* register *) pwire FA_cout_3193;
  (* register *) pwire FA_cout_3194;
  (* register *) pwire FA_cout_3195;
  (* register *) pwire FA_cout_3196;
  (* register *) pwire FA_cout_3197;
  (* register *) pwire FA_cout_3198;
  (* register *) pwire FA_cout_3199;
  (* register *) pwire FA_cout_3200;
  (* register *) pwire FA_cout_3201;
  (* register *) pwire FA_cout_3202;
  (* register *) pwire FA_cout_3203;
  (* register *) pwire FA_cout_3204;
  (* register *) pwire FA_cout_3205;
  (* register *) pwire FA_cout_3206;
  (* register *) pwire FA_cout_3207;
  (* register *) pwire FA_cout_3208;
  (* register *) pwire FA_cout_3209;
  (* register *) pwire FA_cout_3210;
  (* register *) pwire FA_cout_3211;
  (* register *) pwire FA_cout_3212;
  (* register *) pwire FA_cout_3213;
  (* register *) pwire FA_cout_3214;
  (* register *) pwire FA_cout_3215;
  (* register *) pwire FA_cout_3216;
  (* register *) pwire FA_cout_3217;
  (* register *) pwire FA_cout_3218;
  (* register *) pwire FA_cout_3219;
  (* register *) pwire FA_cout_3220;
  (* register *) pwire FA_cout_3221;
  (* register *) pwire FA_cout_3222;
  (* register *) pwire FA_cout_3223;
  (* register *) pwire FA_cout_3224;
  (* register *) pwire FA_cout_3225;
  (* register *) pwire FA_cout_3226;
  (* register *) pwire FA_cout_3227;
  (* register *) pwire FA_cout_3228;
  (* register *) pwire FA_cout_3229;
  (* register *) pwire FA_cout_3230;
  (* register *) pwire FA_cout_3231;
  (* register *) pwire FA_cout_3232;
  (* register *) pwire FA_cout_3233;
  (* register *) pwire FA_cout_3234;
  (* register *) pwire FA_cout_3235;
  (* register *) pwire FA_cout_3236;
  (* register *) pwire FA_cout_3237;
  (* register *) pwire FA_cout_3238;
  (* register *) pwire FA_cout_3239;
  (* register *) pwire FA_cout_3240;
  (* register *) pwire FA_cout_3241;
  (* register *) pwire FA_cout_3242;
  (* register *) pwire FA_cout_3243;
  (* register *) pwire FA_cout_3244;
  (* register *) pwire FA_cout_3245;
  (* register *) pwire FA_cout_3246;
  (* register *) pwire FA_cout_3247;
  (* register *) pwire FA_cout_3248;
  (* register *) pwire FA_cout_3249;
  (* register *) pwire FA_cout_3250;
  (* register *) pwire FA_cout_3251;
  (* register *) pwire FA_cout_3252;
  (* register *) pwire FA_cout_3253;
  (* register *) pwire FA_cout_3254;
  (* register *) pwire FA_cout_3255;
  (* register *) pwire FA_cout_3256;
  (* register *) pwire FA_cout_3257;
  (* register *) pwire FA_cout_3258;
  (* register *) pwire FA_cout_3259;
  (* register *) pwire FA_cout_3260;
  (* register *) pwire FA_cout_3261;
  (* register *) pwire FA_cout_3262;
  (* register *) pwire FA_cout_3263;
  (* register *) pwire FA_cout_3264;
  (* register *) pwire FA_cout_3265;
  (* register *) pwire FA_cout_3266;
  (* register *) pwire FA_cout_3267;
  (* register *) pwire FA_cout_3268;
  (* register *) pwire FA_cout_3269;
  (* register *) pwire FA_cout_3270;
  (* register *) pwire FA_cout_3271;
  (* register *) pwire FA_cout_3272;
  (* register *) pwire FA_cout_3273;
  (* register *) pwire FA_cout_3274;
  (* register *) pwire FA_cout_3275;
  (* register *) pwire FA_cout_3276;
  (* register *) pwire FA_cout_3277;
  (* register *) pwire FA_cout_3278;
  (* register *) pwire FA_cout_3279;
  (* register *) pwire FA_cout_3280;
  (* register *) pwire FA_cout_3281;
  (* register *) pwire FA_cout_3282;
  (* register *) pwire FA_cout_3283;
  (* register *) pwire FA_cout_3284;
  (* register *) pwire FA_cout_3285;
  (* register *) pwire FA_cout_3286;
  (* register *) pwire FA_cout_3287;
  (* register *) pwire FA_cout_3288;
  (* register *) pwire FA_cout_3289;
  (* register *) pwire FA_cout_3290;
  (* register *) pwire FA_cout_3291;
  (* register *) pwire FA_cout_3292;
  (* register *) pwire FA_cout_3293;
  (* register *) pwire FA_cout_3294;
  (* register *) pwire FA_cout_3295;
  (* register *) pwire FA_cout_3296;
  (* register *) pwire FA_cout_3297;
  (* register *) pwire FA_cout_3298;
  (* register *) pwire FA_cout_3299;
  (* register *) pwire FA_cout_3300;
  (* register *) pwire FA_cout_3301;
  (* register *) pwire FA_cout_3302;
  (* register *) pwire FA_cout_3303;
  (* register *) pwire FA_cout_3304;
  (* register *) pwire FA_cout_3305;
  (* register *) pwire FA_cout_3306;
  (* register *) pwire FA_cout_3307;
  (* register *) pwire FA_cout_3308;
  (* register *) pwire FA_cout_3309;
  (* register *) pwire FA_cout_3310;
  (* register *) pwire FA_cout_3311;
  (* register *) pwire FA_cout_3312;
  (* register *) pwire FA_cout_3313;
  (* register *) pwire FA_cout_3314;
  (* register *) pwire FA_cout_3315;
  (* register *) pwire FA_cout_3316;
  (* register *) pwire FA_cout_3317;
  (* register *) pwire FA_cout_3318;
  (* register *) pwire FA_cout_3319;
  (* register *) pwire FA_cout_3320;
  (* register *) pwire FA_cout_3321;
  (* register *) pwire FA_cout_3322;
  (* register *) pwire FA_cout_3323;
  (* register *) pwire FA_cout_3324;
  (* register *) pwire FA_cout_3325;
  (* register *) pwire FA_cout_3326;
  (* register *) pwire FA_cout_3327;
  (* register *) pwire FA_cout_3328;
  (* register *) pwire FA_cout_3329;
  (* register *) pwire FA_cout_3330;
  (* register *) pwire FA_cout_3331;
  (* register *) pwire FA_cout_3332;
  (* register *) pwire FA_cout_3333;
  (* register *) pwire FA_cout_3334;
  (* register *) pwire FA_cout_3335;
  (* register *) pwire FA_cout_3336;
  (* register *) pwire FA_cout_3337;
  (* register *) pwire FA_cout_3338;
  (* register *) pwire FA_cout_3339;
  (* register *) pwire FA_cout_3340;
  (* register *) pwire FA_cout_3341;
  (* register *) pwire FA_cout_3342;
  (* register *) pwire FA_cout_3343;
  (* register *) pwire FA_cout_3344;
  (* register *) pwire FA_cout_3345;
  (* register *) pwire FA_cout_3346;
  (* register *) pwire FA_cout_3347;
  (* register *) pwire FA_cout_3348;
  (* register *) pwire FA_cout_3349;
  (* register *) pwire FA_cout_3350;
  (* register *) pwire FA_cout_3351;
  (* register *) pwire FA_cout_3352;
  (* register *) pwire FA_cout_3353;
  (* register *) pwire FA_cout_3354;
  (* register *) pwire FA_cout_3355;
  (* register *) pwire FA_cout_3356;
  (* register *) pwire FA_cout_3357;
  (* register *) pwire FA_cout_3358;
  (* register *) pwire FA_cout_3359;
  (* register *) pwire FA_cout_3360;
  (* register *) pwire FA_cout_3361;
  (* register *) pwire FA_cout_3362;
  (* register *) pwire FA_cout_3363;
  (* register *) pwire FA_cout_3364;
  (* register *) pwire FA_cout_3365;
  (* register *) pwire FA_cout_3366;
  (* register *) pwire FA_cout_3367;
  (* register *) pwire FA_cout_3368;
  (* register *) pwire FA_cout_3369;
  (* register *) pwire FA_cout_3370;
  (* register *) pwire FA_cout_3371;
  (* register *) pwire FA_cout_3372;
  (* register *) pwire FA_cout_3373;
  (* register *) pwire FA_cout_3374;
  (* register *) pwire FA_cout_3375;
  (* register *) pwire FA_cout_3376;
  (* register *) pwire FA_cout_3377;
  (* register *) pwire FA_cout_3378;
  (* register *) pwire FA_cout_3379;
  (* register *) pwire FA_cout_3380;
  (* register *) pwire FA_cout_3381;
  (* register *) pwire FA_cout_3382;
  (* register *) pwire FA_cout_3383;
  (* register *) pwire FA_cout_3384;
  (* register *) pwire FA_cout_3385;
  (* register *) pwire FA_cout_3386;
  (* register *) pwire FA_cout_3387;
  (* register *) pwire FA_cout_3388;
  (* register *) pwire FA_cout_3389;
  (* register *) pwire FA_cout_3390;
  (* register *) pwire FA_cout_3391;
  (* register *) pwire FA_cout_3392;
  (* register *) pwire FA_cout_3393;
  (* register *) pwire FA_cout_3394;
  (* register *) pwire FA_cout_3395;
  (* register *) pwire FA_cout_3396;
  (* register *) pwire FA_cout_3397;
  (* register *) pwire FA_cout_3398;
  (* register *) pwire FA_cout_3399;
  (* register *) pwire FA_cout_3400;
  (* register *) pwire FA_cout_3401;
  (* register *) pwire FA_cout_3402;
  (* register *) pwire FA_cout_3403;
  (* register *) pwire FA_cout_3404;
  (* register *) pwire FA_cout_3405;
  (* register *) pwire FA_cout_3406;
  (* register *) pwire FA_cout_3407;
  (* register *) pwire FA_cout_3408;
  (* register *) pwire FA_cout_3409;
  (* register *) pwire FA_cout_3410;
  (* register *) pwire FA_cout_3411;
  (* register *) pwire FA_cout_3412;
  (* register *) pwire FA_cout_3413;
  (* register *) pwire FA_cout_3414;
  (* register *) pwire FA_cout_3415;
  (* register *) pwire FA_cout_3416;
  (* register *) pwire FA_cout_3417;
  (* register *) pwire FA_cout_3418;
  (* register *) pwire FA_cout_3419;
  (* register *) pwire FA_cout_3420;
  (* register *) pwire FA_cout_3421;
  (* register *) pwire FA_cout_3422;
  (* register *) pwire FA_cout_3423;
  (* register *) pwire FA_cout_3424;
  (* register *) pwire FA_cout_3425;
  (* register *) pwire FA_cout_3426;
  (* register *) pwire FA_cout_3427;
  (* register *) pwire FA_cout_3428;
  (* register *) pwire FA_cout_3429;
  (* register *) pwire FA_cout_3430;
  (* register *) pwire FA_cout_3431;
  (* register *) pwire FA_cout_3432;
  (* register *) pwire FA_cout_3433;
  (* register *) pwire FA_cout_3434;
  (* register *) pwire FA_cout_3435;
  (* register *) pwire FA_cout_3436;
  (* register *) pwire FA_cout_3437;
  (* register *) pwire FA_cout_3438;
  (* register *) pwire FA_cout_3439;
  (* register *) pwire FA_cout_3440;
  (* register *) pwire FA_cout_3441;
  (* register *) pwire FA_cout_3442;
  (* register *) pwire FA_cout_3443;
  (* register *) pwire FA_cout_3444;
  (* register *) pwire FA_cout_3445;
  (* register *) pwire FA_cout_3446;
  (* register *) pwire FA_cout_3447;
  (* register *) pwire FA_cout_3448;
  (* register *) pwire FA_cout_3449;
  (* register *) pwire FA_cout_3450;
  (* register *) pwire FA_cout_3451;
  (* register *) pwire FA_cout_3452;
  (* register *) pwire FA_cout_3453;
  (* register *) pwire FA_cout_3454;
  (* register *) pwire FA_cout_3455;
  (* register *) pwire FA_cout_3456;
  (* register *) pwire FA_cout_3457;
  (* register *) pwire FA_cout_3458;
  (* register *) pwire FA_cout_3459;
  (* register *) pwire FA_cout_3460;
  (* register *) pwire FA_cout_3461;
  (* register *) pwire FA_cout_3462;
  (* register *) pwire FA_cout_3463;
  (* register *) pwire FA_cout_3464;
  (* register *) pwire FA_cout_3465;
  (* register *) pwire FA_cout_3466;
  (* register *) pwire FA_cout_3467;
  (* register *) pwire FA_cout_3468;
  (* register *) pwire FA_cout_3469;
  (* register *) pwire FA_cout_3470;
  (* register *) pwire FA_cout_3471;
  (* register *) pwire FA_cout_3472;
  (* register *) pwire FA_cout_3473;
  (* register *) pwire FA_cout_3474;
  (* register *) pwire FA_cout_3475;
  (* register *) pwire FA_cout_3476;
  (* register *) pwire FA_cout_3477;
  (* register *) pwire FA_cout_3478;
  (* register *) pwire FA_cout_3479;
  (* register *) pwire FA_cout_3480;
  (* register *) pwire FA_cout_3481;
  (* register *) pwire FA_cout_3482;
  (* register *) pwire FA_cout_3483;
  (* register *) pwire FA_cout_3484;
  (* register *) pwire FA_cout_3485;
  (* register *) pwire FA_cout_3486;
  (* register *) pwire FA_cout_3487;
  (* register *) pwire FA_cout_3488;
  (* register *) pwire FA_cout_3489;
  (* register *) pwire FA_cout_3490;
  (* register *) pwire FA_cout_3491;
  (* register *) pwire FA_cout_3492;
  (* register *) pwire FA_cout_3493;
  (* register *) pwire FA_cout_3494;
  (* register *) pwire FA_cout_3495;
  (* register *) pwire FA_cout_3496;
  (* register *) pwire FA_cout_3497;
  (* register *) pwire FA_cout_3498;
  (* register *) pwire FA_cout_3499;
  (* register *) pwire FA_cout_3500;
  (* register *) pwire FA_cout_3501;
  (* register *) pwire FA_cout_3502;
  (* register *) pwire FA_cout_3503;
  (* register *) pwire FA_cout_3504;
  (* register *) pwire FA_cout_3505;
  (* register *) pwire FA_cout_3506;
  (* register *) pwire FA_cout_3507;
  (* register *) pwire FA_cout_3508;
  (* register *) pwire FA_cout_3509;
  (* register *) pwire FA_cout_3510;
  (* register *) pwire FA_cout_3511;
  (* register *) pwire FA_cout_3512;
  (* register *) pwire FA_cout_3513;
  (* register *) pwire FA_cout_3514;
  (* register *) pwire FA_cout_3515;
  (* register *) pwire FA_cout_3516;
  (* register *) pwire FA_cout_3517;
  (* register *) pwire FA_cout_3518;
  (* register *) pwire FA_cout_3519;
  (* register *) pwire FA_cout_3520;
  (* register *) pwire FA_cout_3521;
  (* register *) pwire FA_cout_3522;
  (* register *) pwire FA_cout_3523;
  (* register *) pwire FA_cout_3524;
  (* register *) pwire FA_cout_3525;
  (* register *) pwire FA_cout_3526;
  (* register *) pwire FA_cout_3527;
  (* register *) pwire FA_cout_3528;
  (* register *) pwire FA_cout_3529;
  (* register *) pwire FA_cout_3530;
  (* register *) pwire FA_cout_3531;
  (* register *) pwire FA_cout_3532;
  (* register *) pwire FA_cout_3533;
  (* register *) pwire FA_cout_3534;
  (* register *) pwire FA_cout_3535;
  (* register *) pwire FA_cout_3536;
  (* register *) pwire FA_cout_3537;
  (* register *) pwire FA_cout_3538;
  (* register *) pwire FA_cout_3539;
  (* register *) pwire FA_cout_3540;
  (* register *) pwire FA_cout_3541;
  (* register *) pwire FA_cout_3542;
  (* register *) pwire FA_cout_3543;
  (* register *) pwire FA_cout_3544;
  (* register *) pwire FA_cout_3545;
  (* register *) pwire FA_cout_3546;
  (* register *) pwire FA_cout_3547;
  (* register *) pwire FA_cout_3548;
  (* register *) pwire FA_cout_3549;
  (* register *) pwire FA_cout_3550;
  (* register *) pwire FA_cout_3551;
  (* register *) pwire FA_cout_3552;
  (* register *) pwire FA_cout_3553;
  (* register *) pwire FA_cout_3554;
  (* register *) pwire FA_cout_3555;
  (* register *) pwire FA_cout_3556;
  (* register *) pwire FA_cout_3557;
  (* register *) pwire FA_cout_3558;
  (* register *) pwire FA_cout_3559;
  (* register *) pwire FA_cout_3560;
  (* register *) pwire FA_cout_3561;
  (* register *) pwire FA_cout_3562;
  (* register *) pwire FA_cout_3563;
  (* register *) pwire FA_cout_3564;
  (* register *) pwire FA_cout_3565;
  (* register *) pwire FA_cout_3566;
  (* register *) pwire FA_cout_3567;
  (* register *) pwire FA_cout_3568;
  (* register *) pwire FA_cout_3569;
  (* register *) pwire FA_cout_3570;
  (* register *) pwire FA_cout_3571;
  (* register *) pwire FA_cout_3572;
  (* register *) pwire FA_cout_3573;
  (* register *) pwire FA_cout_3574;
  (* register *) pwire FA_cout_3575;
  (* register *) pwire FA_cout_3576;
  (* register *) pwire FA_cout_3577;
  (* register *) pwire FA_cout_3578;
  (* register *) pwire FA_cout_3579;
  (* register *) pwire FA_cout_3580;
  (* register *) pwire FA_cout_3581;
  (* register *) pwire FA_cout_3582;
  (* register *) pwire FA_cout_3583;
  (* register *) pwire FA_cout_3584;
  (* register *) pwire FA_cout_3585;
  (* register *) pwire FA_cout_3586;
  (* register *) pwire FA_cout_3587;
  (* register *) pwire FA_cout_3588;
  (* register *) pwire FA_cout_3589;
  (* register *) pwire FA_cout_3590;
  (* register *) pwire FA_cout_3591;
  (* register *) pwire FA_cout_3592;
  (* register *) pwire FA_cout_3593;
  (* register *) pwire FA_cout_3594;
  (* register *) pwire FA_cout_3595;
  (* register *) pwire FA_cout_3596;
  (* register *) pwire FA_cout_3597;
  (* register *) pwire FA_cout_3598;
  (* register *) pwire FA_cout_3599;
  (* register *) pwire FA_cout_3600;
  (* register *) pwire FA_cout_3601;
  (* register *) pwire FA_cout_3602;
  (* register *) pwire FA_cout_3603;
  (* register *) pwire FA_cout_3604;
  (* register *) pwire FA_cout_3605;
  (* register *) pwire FA_cout_3606;
  (* register *) pwire FA_cout_3607;
  (* register *) pwire FA_cout_3608;
  (* register *) pwire FA_cout_3609;
  (* register *) pwire FA_cout_3610;
  (* register *) pwire FA_cout_3611;
  (* register *) pwire FA_cout_3612;
  (* register *) pwire FA_cout_3613;
  (* register *) pwire FA_cout_3614;
  (* register *) pwire FA_cout_3615;
  (* register *) pwire FA_cout_3616;
  (* register *) pwire FA_cout_3617;
  (* register *) pwire FA_cout_3618;
  (* register *) pwire FA_cout_3619;
  (* register *) pwire FA_cout_3620;
  (* register *) pwire FA_cout_3621;
  (* register *) pwire FA_cout_3622;
  (* register *) pwire FA_cout_3623;
  (* register *) pwire FA_cout_3624;
  (* register *) pwire FA_cout_3625;
  (* register *) pwire FA_cout_3626;
  (* register *) pwire FA_cout_3627;
  (* register *) pwire FA_cout_3628;
  (* register *) pwire FA_cout_3629;
  (* register *) pwire FA_cout_3630;
  (* register *) pwire FA_cout_3631;
  (* register *) pwire FA_cout_3632;
  (* register *) pwire FA_cout_3633;
  (* register *) pwire FA_cout_3634;
  (* register *) pwire FA_cout_3635;
  (* register *) pwire FA_cout_3636;
  (* register *) pwire FA_cout_3637;
  (* register *) pwire FA_cout_3638;
  (* register *) pwire FA_cout_3639;
  (* register *) pwire FA_cout_3640;
  (* register *) pwire FA_cout_3641;
  (* register *) pwire FA_cout_3642;
  (* register *) pwire FA_cout_3643;
  (* register *) pwire FA_cout_3644;
  (* register *) pwire FA_cout_3645;
  (* register *) pwire FA_cout_3646;
  (* register *) pwire FA_cout_3647;
  (* register *) pwire FA_cout_3648;
  (* register *) pwire FA_cout_3649;
  (* register *) pwire FA_cout_3650;
  (* register *) pwire FA_cout_3651;
  (* register *) pwire FA_cout_3652;
  (* register *) pwire FA_cout_3653;
  (* register *) pwire FA_cout_3654;
  (* register *) pwire FA_cout_3655;
  (* register *) pwire FA_cout_3656;
  (* register *) pwire FA_cout_3657;
  (* register *) pwire FA_cout_3658;
  (* register *) pwire FA_cout_3659;
  (* register *) pwire FA_cout_3660;
  (* register *) pwire FA_cout_3661;
  (* register *) pwire FA_cout_3662;
  (* register *) pwire FA_cout_3663;
  (* register *) pwire FA_cout_3664;
  (* register *) pwire FA_cout_3665;
  (* register *) pwire FA_cout_3666;
  (* register *) pwire FA_cout_3667;
  (* register *) pwire FA_cout_3668;
  (* register *) pwire FA_cout_3669;
  (* register *) pwire FA_cout_3670;
  (* register *) pwire FA_cout_3671;
  (* register *) pwire FA_cout_3672;
  (* register *) pwire FA_cout_3673;
  (* register *) pwire FA_cout_3674;
  (* register *) pwire FA_cout_3675;
  (* register *) pwire FA_cout_3676;
  (* register *) pwire FA_cout_3677;
  (* register *) pwire FA_cout_3678;
  (* register *) pwire FA_cout_3679;
  (* register *) pwire FA_cout_3680;
  (* register *) pwire FA_cout_3681;
  (* register *) pwire FA_cout_3682;
  (* register *) pwire FA_cout_3683;
  (* register *) pwire FA_cout_3684;
  (* register *) pwire FA_cout_3685;
  (* register *) pwire FA_cout_3686;
  (* register *) pwire FA_cout_3687;
  (* register *) pwire FA_cout_3688;
  (* register *) pwire FA_cout_3689;
  (* register *) pwire FA_cout_3690;
  (* register *) pwire FA_cout_3691;
  (* register *) pwire FA_cout_3692;
  (* register *) pwire FA_cout_3693;
  (* register *) pwire FA_cout_3694;
  (* register *) pwire FA_cout_3695;
  (* register *) pwire FA_cout_3696;
  (* register *) pwire FA_cout_3697;
  (* register *) pwire FA_cout_3698;
  (* register *) pwire FA_cout_3699;
  (* register *) pwire FA_cout_3700;
  (* register *) pwire FA_cout_3701;
  (* register *) pwire FA_cout_3702;
  (* register *) pwire FA_cout_3703;
  (* register *) pwire FA_cout_3704;
  (* register *) pwire FA_cout_3705;
  (* register *) pwire FA_cout_3706;
  (* register *) pwire FA_cout_3707;
  (* register *) pwire FA_cout_3708;
  (* register *) pwire FA_cout_3709;
  (* register *) pwire FA_cout_3710;
  (* register *) pwire FA_cout_3711;
  (* register *) pwire FA_cout_3712;
  (* register *) pwire FA_cout_3713;
  (* register *) pwire FA_cout_3714;
  (* register *) pwire FA_cout_3715;
  (* register *) pwire FA_cout_3716;
  (* register *) pwire FA_cout_3717;
  (* register *) pwire FA_cout_3718;
  (* register *) pwire FA_cout_3719;
  (* register *) pwire FA_cout_3720;
  (* register *) pwire FA_cout_3721;
  (* register *) pwire FA_cout_3722;
  (* register *) pwire FA_cout_3723;
  (* register *) pwire FA_cout_3724;
  (* register *) pwire FA_cout_3725;
  (* register *) pwire FA_cout_3726;
  (* register *) pwire FA_cout_3727;
  (* register *) pwire FA_cout_3728;
  (* register *) pwire FA_cout_3729;
  (* register *) pwire FA_cout_3730;
  (* register *) pwire FA_cout_3731;
  (* register *) pwire FA_cout_3732;
  (* register *) pwire FA_cout_3733;
  (* register *) pwire FA_cout_3734;
  (* register *) pwire FA_cout_3735;
  (* register *) pwire FA_cout_3736;
  (* register *) pwire FA_cout_3737;
  (* register *) pwire FA_cout_3738;
  (* register *) pwire FA_cout_3739;
  (* register *) pwire FA_cout_3740;
  (* register *) pwire FA_cout_3741;
  (* register *) pwire FA_cout_3742;
  (* register *) pwire FA_cout_3743;
  (* register *) pwire FA_cout_3744;
  (* register *) pwire FA_cout_3745;
  (* register *) pwire FA_cout_3746;
  (* register *) pwire FA_cout_3747;
  (* register *) pwire FA_cout_3748;
  (* register *) pwire FA_cout_3749;
  (* register *) pwire FA_cout_3750;
  (* register *) pwire FA_cout_3751;
  (* register *) pwire FA_cout_3752;
  (* register *) pwire FA_cout_3753;
  (* register *) pwire FA_cout_3754;
  (* register *) pwire FA_cout_3755;
  (* register *) pwire FA_cout_3756;
  (* register *) pwire FA_cout_3757;
  (* register *) pwire FA_cout_3758;
  (* register *) pwire FA_cout_3759;
  (* register *) pwire FA_cout_3760;
  (* register *) pwire FA_cout_3761;
  (* register *) pwire FA_cout_3762;
  (* register *) pwire FA_cout_3763;
  (* register *) pwire FA_cout_3764;
  (* register *) pwire FA_cout_3765;
  (* register *) pwire FA_cout_3766;
  (* register *) pwire FA_cout_3767;
  (* register *) pwire FA_cout_3768;
  (* register *) pwire FA_cout_3769;
  (* register *) pwire FA_cout_3770;
  (* register *) pwire FA_cout_3771;
  (* register *) pwire FA_cout_3772;
  (* register *) pwire FA_cout_3773;
  (* register *) pwire FA_cout_3774;
  (* register *) pwire FA_cout_3775;
  (* register *) pwire FA_cout_3776;
  (* register *) pwire FA_cout_3777;
  (* register *) pwire FA_cout_3778;
  (* register *) pwire FA_cout_3779;
  (* register *) pwire FA_cout_3780;
  (* register *) pwire FA_cout_3781;
  (* register *) pwire FA_cout_3782;
  (* register *) pwire FA_cout_3783;
  (* register *) pwire FA_cout_3784;
  (* register *) pwire FA_cout_3785;
  (* register *) pwire FA_cout_3786;
  (* register *) pwire FA_cout_3787;
  (* register *) pwire FA_cout_3788;
  (* register *) pwire FA_cout_3789;
  (* register *) pwire FA_cout_3790;
  (* register *) pwire FA_cout_3791;
  (* register *) pwire FA_cout_3792;
  (* register *) pwire FA_cout_3793;
  (* register *) pwire FA_cout_3794;
  (* register *) pwire FA_cout_3795;
  (* register *) pwire FA_cout_3796;
  (* register *) pwire FA_cout_3797;
  (* register *) pwire FA_cout_3798;
  (* register *) pwire FA_cout_3799;
  (* register *) pwire FA_cout_3800;
  (* register *) pwire FA_cout_3801;
  (* register *) pwire FA_cout_3802;
  (* register *) pwire FA_cout_3803;
  (* register *) pwire FA_cout_3804;
  (* register *) pwire FA_cout_3805;
  (* register *) pwire FA_cout_3806;
  (* register *) pwire FA_cout_3807;
  (* register *) pwire FA_cout_3808;
  (* register *) pwire FA_cout_3809;
  (* register *) pwire FA_cout_3810;
  (* register *) pwire FA_cout_3811;
  (* register *) pwire FA_cout_3812;
  (* register *) pwire FA_cout_3813;
  (* register *) pwire FA_cout_3814;
  (* register *) pwire FA_cout_3815;
  (* register *) pwire FA_cout_3816;
  (* register *) pwire FA_cout_3817;
  (* register *) pwire FA_cout_3818;
  (* register *) pwire FA_cout_3819;
  (* register *) pwire FA_cout_3820;
  (* register *) pwire FA_cout_3821;
  (* register *) pwire FA_cout_3822;
  (* register *) pwire FA_cout_3823;
  (* register *) pwire FA_cout_3824;
  (* register *) pwire FA_cout_3825;
  (* register *) pwire FA_cout_3826;
  (* register *) pwire FA_cout_3827;
  (* register *) pwire FA_cout_3828;
  (* register *) pwire FA_cout_3829;
  (* register *) pwire FA_cout_3830;
  (* register *) pwire FA_cout_3831;
  (* register *) pwire FA_cout_3832;
  (* register *) pwire FA_cout_3833;
  (* register *) pwire FA_cout_3834;
  (* register *) pwire FA_cout_3835;
  (* register *) pwire FA_cout_3836;
  (* register *) pwire FA_cout_3837;
  (* register *) pwire FA_cout_3838;
  (* register *) pwire FA_cout_3839;
  (* register *) pwire FA_cout_3840;
  (* register *) pwire FA_cout_3841;
  (* register *) pwire FA_cout_3842;
  (* register *) pwire FA_cout_3843;
  (* register *) pwire FA_cout_3844;
  (* register *) pwire FA_cout_3845;
  (* register *) pwire HA_out_0;
  (* register *) pwire HA_out_1;
  (* register *) pwire HA_out_2;
  (* register *) pwire HA_out_3;
  (* register *) pwire HA_out_4;
  (* register *) pwire HA_out_5;
  (* register *) pwire HA_out_6;
  (* register *) pwire HA_out_7;
  (* register *) pwire HA_out_8;
  (* register *) pwire HA_out_9;
  (* register *) pwire HA_out_10;
  (* register *) pwire HA_out_11;
  (* register *) pwire HA_out_12;
  (* register *) pwire HA_out_13;
  (* register *) pwire HA_out_14;
  (* register *) pwire HA_out_15;
  (* register *) pwire HA_out_16;
  (* register *) pwire HA_out_17;
  (* register *) pwire HA_out_18;
  (* register *) pwire HA_out_19;
  (* register *) pwire HA_out_20;
  (* register *) pwire HA_out_21;
  (* register *) pwire HA_out_22;
  (* register *) pwire HA_out_23;
  (* register *) pwire HA_out_24;
  (* register *) pwire HA_out_25;
  (* register *) pwire HA_out_26;
  (* register *) pwire HA_out_27;
  (* register *) pwire HA_out_28;
  (* register *) pwire HA_out_29;
  (* register *) pwire HA_out_30;
  (* register *) pwire HA_out_31;
  (* register *) pwire HA_out_32;
  (* register *) pwire HA_out_33;
  (* register *) pwire HA_out_34;
  (* register *) pwire HA_out_35;
  (* register *) pwire HA_out_36;
  (* register *) pwire HA_out_37;
  (* register *) pwire HA_out_38;
  (* register *) pwire HA_out_39;
  (* register *) pwire HA_out_40;
  (* register *) pwire HA_out_41;
  (* register *) pwire HA_out_42;
  (* register *) pwire HA_out_43;
  (* register *) pwire HA_out_44;
  (* register *) pwire HA_out_45;
  (* register *) pwire HA_out_46;
  (* register *) pwire HA_out_47;
  (* register *) pwire HA_out_48;
  (* register *) pwire HA_out_49;
  (* register *) pwire HA_out_50;
  (* register *) pwire HA_out_51;
  (* register *) pwire HA_out_52;
  (* register *) pwire HA_out_53;
  (* register *) pwire HA_out_54;
  (* register *) pwire HA_out_55;
  (* register *) pwire HA_out_56;
  (* register *) pwire HA_out_57;
  (* register *) pwire HA_out_58;
  (* register *) pwire HA_out_59;
  (* register *) pwire HA_out_60;
  (* register *) pwire HA_out_61;
  (* register *) pwire HA_out_62;
  (* register *) pwire HA_out_63;
  (* register *) pwire HA_out_64;
  (* register *) pwire HA_out_65;
  (* register *) pwire HA_out_66;
  (* register *) pwire HA_out_67;
  (* register *) pwire HA_out_68;
  (* register *) pwire HA_out_69;
  (* register *) pwire HA_out_70;
  (* register *) pwire HA_out_71;
  (* register *) pwire HA_out_72;
  (* register *) pwire HA_out_73;
  (* register *) pwire HA_out_74;
  (* register *) pwire HA_out_75;
  (* register *) pwire HA_out_76;
  (* register *) pwire HA_out_77;
  (* register *) pwire HA_out_78;
  (* register *) pwire HA_out_79;
  (* register *) pwire HA_out_80;
  (* register *) pwire HA_out_81;
  (* register *) pwire HA_out_82;
  (* register *) pwire HA_out_83;
  (* register *) pwire HA_out_84;
  (* register *) pwire HA_out_85;
  (* register *) pwire HA_out_86;
  (* register *) pwire HA_out_87;
  (* register *) pwire HA_out_88;
  (* register *) pwire HA_out_89;
  (* register *) pwire HA_out_90;
  (* register *) pwire HA_out_91;
  (* register *) pwire HA_out_92;
  (* register *) pwire HA_out_93;
  (* register *) pwire HA_out_94;
  (* register *) pwire HA_out_95;
  (* register *) pwire HA_out_96;
  (* register *) pwire HA_out_97;
  (* register *) pwire HA_out_98;
  (* register *) pwire HA_out_99;
  (* register *) pwire HA_out_100;
  (* register *) pwire HA_out_101;
  (* register *) pwire HA_out_102;
  (* register *) pwire HA_out_103;
  (* register *) pwire HA_out_104;
  (* register *) pwire HA_out_105;
  (* register *) pwire HA_out_106;
  (* register *) pwire HA_out_107;
  (* register *) pwire HA_out_108;
  (* register *) pwire HA_out_109;
  (* register *) pwire HA_out_110;
  (* register *) pwire HA_out_111;
  (* register *) pwire HA_out_112;
  (* register *) pwire HA_out_113;
  (* register *) pwire HA_out_114;
  (* register *) pwire HA_out_115;
  (* register *) pwire HA_out_116;
  (* register *) pwire HA_out_117;
  (* register *) pwire HA_out_118;
  (* register *) pwire HA_out_119;
  (* register *) pwire HA_out_120;
  (* register *) pwire HA_out_121;
  (* register *) pwire HA_out_122;
  (* register *) pwire HA_out_123;
  (* register *) pwire HA_out_124;
  (* register *) pwire HA_out_125;
  (* register *) pwire HA_out_126;
  (* register *) pwire HA_out_127;
  (* register *) pwire HA_out_128;
  (* register *) pwire HA_out_129;
  (* register *) pwire HA_out_130;
  (* register *) pwire HA_out_131;
  (* register *) pwire HA_out_132;
  (* register *) pwire HA_out_133;
  (* register *) pwire HA_out_134;
  (* register *) pwire HA_out_135;
  (* register *) pwire HA_out_136;
  (* register *) pwire HA_out_137;
  (* register *) pwire HA_out_138;
  (* register *) pwire HA_out_139;
  (* register *) pwire HA_out_140;
  (* register *) pwire HA_out_141;
  (* register *) pwire HA_out_142;
  (* register *) pwire HA_out_143;
  (* register *) pwire HA_out_144;
  (* register *) pwire HA_out_145;
  (* register *) pwire HA_out_146;
  (* register *) pwire HA_out_147;
  (* register *) pwire HA_out_148;
  (* register *) pwire HA_out_149;
  (* register *) pwire HA_out_150;
  (* register *) pwire HA_out_151;
  (* register *) pwire HA_out_152;
  (* register *) pwire HA_out_153;
  (* register *) pwire HA_out_154;
  (* register *) pwire HA_out_155;
  (* register *) pwire HA_out_156;
  (* register *) pwire HA_out_157;
  (* register *) pwire HA_out_158;
  (* register *) pwire HA_out_159;
  (* register *) pwire HA_out_160;
  (* register *) pwire HA_out_161;
  (* register *) pwire HA_out_162;
  (* register *) pwire HA_out_163;
  (* register *) pwire HA_out_164;
  (* register *) pwire HA_out_165;
  (* register *) pwire HA_out_166;
  (* register *) pwire HA_out_167;
  (* register *) pwire HA_out_168;
  (* register *) pwire HA_out_169;
  (* register *) pwire HA_out_170;
  (* register *) pwire HA_out_171;
  (* register *) pwire HA_out_172;
  (* register *) pwire HA_out_173;
  (* register *) pwire HA_out_174;
  (* register *) pwire HA_out_175;
  (* register *) pwire HA_out_176;
  (* register *) pwire HA_out_177;
  (* register *) pwire HA_out_178;
  (* register *) pwire HA_out_179;
  (* register *) pwire HA_out_180;
  (* register *) pwire HA_out_181;
  (* register *) pwire HA_out_182;
  (* register *) pwire HA_out_183;
  (* register *) pwire HA_out_184;
  (* register *) pwire HA_out_185;
  (* register *) pwire HA_out_186;
  (* register *) pwire HA_out_187;
  (* register *) pwire HA_out_188;
  (* register *) pwire HA_out_189;
  (* register *) pwire HA_out_190;
  (* register *) pwire HA_out_191;
  (* register *) pwire HA_out_192;
  (* register *) pwire HA_out_193;
  (* register *) pwire HA_out_194;
  (* register *) pwire HA_out_195;
  (* register *) pwire HA_out_196;
  (* register *) pwire HA_out_197;
  (* register *) pwire HA_out_198;
  (* register *) pwire HA_out_199;
  (* register *) pwire HA_out_200;
  (* register *) pwire HA_out_201;
  (* register *) pwire HA_out_202;
  (* register *) pwire HA_out_203;
  (* register *) pwire HA_out_204;
  (* register *) pwire HA_out_205;
  (* register *) pwire HA_out_206;
  (* register *) pwire HA_out_207;
  (* register *) pwire HA_out_208;
  (* register *) pwire HA_out_209;
  (* register *) pwire HA_out_210;
  (* register *) pwire HA_out_211;
  (* register *) pwire HA_out_212;
  (* register *) pwire HA_out_213;
  (* register *) pwire HA_out_214;
  (* register *) pwire HA_out_215;
  (* register *) pwire HA_out_216;
  (* register *) pwire HA_out_217;
  (* register *) pwire HA_out_218;
  (* register *) pwire HA_out_219;
  (* register *) pwire HA_out_220;
  (* register *) pwire HA_out_221;
  (* register *) pwire HA_out_222;
  (* register *) pwire HA_out_223;
  (* register *) pwire HA_out_224;
  (* register *) pwire HA_out_225;
  (* register *) pwire HA_out_226;
  (* register *) pwire HA_out_227;
  (* register *) pwire HA_out_228;
  (* register *) pwire HA_out_229;
  (* register *) pwire HA_out_230;
  (* register *) pwire HA_out_231;
  (* register *) pwire HA_out_232;
  (* register *) pwire HA_out_233;
  (* register *) pwire HA_out_234;
  (* register *) pwire HA_out_235;
  (* register *) pwire HA_out_236;
  (* register *) pwire HA_out_237;
  (* register *) pwire HA_out_238;
  (* register *) pwire HA_out_239;
  (* register *) pwire HA_out_240;
  (* register *) pwire HA_out_241;
  (* register *) pwire HA_out_242;
  (* register *) pwire HA_out_243;
  (* register *) pwire HA_out_244;
  (* register *) pwire HA_out_245;
  (* register *) pwire HA_out_246;
  (* register *) pwire HA_out_247;
  (* register *) pwire HA_out_248;
  (* register *) pwire HA_out_249;
  (* register *) pwire HA_out_250;
  (* register *) pwire HA_out_251;
  (* register *) pwire HA_out_252;
  (* register *) pwire HA_out_253;
  (* register *) pwire HA_out_254;
  (* register *) pwire HA_out_255;
  (* register *) pwire HA_out_256;
  (* register *) pwire HA_out_257;
  (* register *) pwire HA_out_258;
  (* register *) pwire HA_out_259;
  (* register *) pwire HA_out_260;
  (* register *) pwire HA_out_261;
  (* register *) pwire HA_out_262;
  (* register *) pwire HA_out_263;
  (* register *) pwire HA_out_264;
  (* register *) pwire HA_out_265;
  (* register *) pwire HA_out_266;
  (* register *) pwire HA_out_267;
  (* register *) pwire HA_out_268;
  (* register *) pwire HA_out_269;
  (* register *) pwire HA_out_270;
  (* register *) pwire HA_out_271;
  (* register *) pwire HA_out_272;
  (* register *) pwire HA_out_273;
  (* register *) pwire HA_out_274;
  (* register *) pwire HA_out_275;
  (* register *) pwire HA_out_276;
  (* register *) pwire HA_out_277;
  (* register *) pwire HA_out_278;
  (* register *) pwire HA_out_279;
  (* register *) pwire HA_out_280;
  (* register *) pwire HA_out_281;
  (* register *) pwire HA_out_282;
  (* register *) pwire HA_out_283;
  (* register *) pwire HA_out_284;
  (* register *) pwire HA_out_285;
  (* register *) pwire HA_out_286;
  (* register *) pwire HA_out_287;
  (* register *) pwire HA_out_288;
  (* register *) pwire HA_out_289;
  (* register *) pwire HA_out_290;
  (* register *) pwire HA_out_291;
  (* register *) pwire HA_out_292;
  (* register *) pwire HA_out_293;
  (* register *) pwire HA_out_294;
  (* register *) pwire HA_out_295;
  (* register *) pwire HA_out_296;
  (* register *) pwire HA_out_297;
  (* register *) pwire HA_out_298;
  (* register *) pwire HA_out_299;
  (* register *) pwire HA_out_300;
  (* register *) pwire HA_out_301;
  (* register *) pwire HA_out_302;
  (* register *) pwire HA_out_303;
  (* register *) pwire HA_out_304;
  (* register *) pwire HA_out_305;
  (* register *) pwire HA_out_306;
  (* register *) pwire HA_out_307;
  (* register *) pwire HA_out_308;
  (* register *) pwire HA_out_309;
  (* register *) pwire HA_out_310;
  (* register *) pwire HA_out_311;
  (* register *) pwire HA_out_312;
  (* register *) pwire HA_out_313;
  (* register *) pwire HA_out_314;
  (* register *) pwire HA_out_315;
  (* register *) pwire HA_out_316;
  (* register *) pwire HA_out_317;
  (* register *) pwire HA_out_318;
  (* register *) pwire HA_out_319;
  (* register *) pwire HA_out_320;
  (* register *) pwire HA_out_321;
  (* register *) pwire HA_out_322;
  (* register *) pwire HA_out_323;
  (* register *) pwire HA_out_324;
  (* register *) pwire HA_out_325;
  (* register *) pwire HA_out_326;
  (* register *) pwire HA_out_327;
  (* register *) pwire HA_out_328;
  (* register *) pwire HA_out_329;
  (* register *) pwire HA_out_330;
  (* register *) pwire HA_out_331;
  (* register *) pwire HA_out_332;
  (* register *) pwire HA_out_333;
  (* register *) pwire HA_out_334;
  (* register *) pwire HA_out_335;
  (* register *) pwire HA_out_336;
  (* register *) pwire HA_out_337;
  (* register *) pwire HA_out_338;
  (* register *) pwire HA_out_339;
  (* register *) pwire HA_out_340;
  (* register *) pwire HA_out_341;
  (* register *) pwire HA_out_342;
  (* register *) pwire HA_out_343;
  (* register *) pwire HA_out_344;
  (* register *) pwire HA_out_345;
  (* register *) pwire HA_out_346;
  (* register *) pwire HA_out_347;
  (* register *) pwire HA_out_348;
  (* register *) pwire HA_out_349;
  (* register *) pwire HA_out_350;
  (* register *) pwire HA_out_351;
  (* register *) pwire HA_out_352;
  (* register *) pwire HA_out_353;
  (* register *) pwire HA_out_354;
  (* register *) pwire HA_out_355;
  (* register *) pwire HA_out_356;
  (* register *) pwire HA_out_357;
  (* register *) pwire HA_out_358;
  (* register *) pwire HA_out_359;
  (* register *) pwire HA_out_360;
  (* register *) pwire HA_out_361;
  (* register *) pwire HA_out_362;
  (* register *) pwire HA_out_363;
  (* register *) pwire HA_out_364;
  (* register *) pwire HA_out_365;
  (* register *) pwire HA_out_366;
  (* register *) pwire HA_out_367;
  (* register *) pwire HA_out_368;
  (* register *) pwire HA_out_369;
  (* register *) pwire HA_out_370;
  (* register *) pwire HA_out_371;
  (* register *) pwire HA_out_372;
  (* register *) pwire HA_out_373;
  (* register *) pwire HA_out_374;
  (* register *) pwire HA_out_375;
  (* register *) pwire HA_out_376;
  (* register *) pwire HA_out_377;
  (* register *) pwire HA_out_378;
  (* register *) pwire HA_out_379;
  (* register *) pwire HA_out_380;
  (* register *) pwire HA_out_381;
  (* register *) pwire HA_out_382;
  (* register *) pwire HA_out_383;
  (* register *) pwire HA_out_384;
  (* register *) pwire HA_out_385;
  (* register *) pwire HA_out_386;
  (* register *) pwire HA_out_387;
  (* register *) pwire HA_out_388;
  (* register *) pwire HA_out_389;
  (* register *) pwire HA_out_390;
  (* register *) pwire HA_out_391;
  (* register *) pwire HA_out_392;
  (* register *) pwire HA_out_393;
  (* register *) pwire HA_out_394;
  (* register *) pwire HA_out_395;
  (* register *) pwire HA_out_396;
  (* register *) pwire HA_out_397;
  (* register *) pwire HA_out_398;
  (* register *) pwire HA_out_399;
  (* register *) pwire HA_out_400;
  (* register *) pwire HA_out_401;
  (* register *) pwire HA_out_402;
  (* register *) pwire HA_out_403;
  (* register *) pwire HA_out_404;
  (* register *) pwire HA_out_405;
  (* register *) pwire HA_out_406;
  (* register *) pwire HA_out_407;
  (* register *) pwire HA_out_408;
  (* register *) pwire HA_out_409;
  (* register *) pwire HA_out_410;
  (* register *) pwire HA_out_411;
  (* register *) pwire HA_out_412;
  (* register *) pwire HA_out_413;
  (* register *) pwire HA_out_414;
  (* register *) pwire HA_out_415;
  (* register *) pwire HA_out_416;
  (* register *) pwire HA_out_417;
  (* register *) pwire HA_out_418;
  (* register *) pwire HA_out_419;
  (* register *) pwire HA_out_420;
  (* register *) pwire HA_out_421;
  (* register *) pwire HA_out_422;
  (* register *) pwire HA_out_423;
  (* register *) pwire HA_out_424;
  (* register *) pwire HA_out_425;
  (* register *) pwire HA_out_426;
  (* register *) pwire HA_out_427;
  (* register *) pwire HA_out_428;
  (* register *) pwire HA_out_429;
  (* register *) pwire HA_out_430;
  (* register *) pwire HA_out_431;
  (* register *) pwire HA_out_432;
  (* register *) pwire HA_out_433;
  (* register *) pwire HA_out_434;
  (* register *) pwire HA_out_435;
  (* register *) pwire HA_out_436;
  (* register *) pwire HA_out_437;
  (* register *) pwire HA_out_438;
  (* register *) pwire HA_out_439;
  (* register *) pwire HA_out_440;
  (* register *) pwire HA_out_441;
  (* register *) pwire HA_out_442;
  (* register *) pwire HA_out_443;
  (* register *) pwire HA_out_444;
  (* register *) pwire HA_out_445;
  (* register *) pwire HA_out_446;
  (* register *) pwire HA_out_447;
  (* register *) pwire HA_out_448;
  (* register *) pwire HA_out_449;
  (* register *) pwire HA_out_450;
  (* register *) pwire HA_out_451;
  (* register *) pwire HA_out_452;
  (* register *) pwire HA_out_453;
  (* register *) pwire HA_out_454;
  (* register *) pwire HA_out_455;
  (* register *) pwire HA_out_456;
  (* register *) pwire HA_out_457;
  (* register *) pwire HA_out_458;
  (* register *) pwire HA_out_459;
  (* register *) pwire HA_out_460;
  (* register *) pwire HA_out_461;
  (* register *) pwire HA_out_462;
  (* register *) pwire HA_out_463;
  (* register *) pwire HA_out_464;
  (* register *) pwire HA_out_465;
  (* register *) pwire HA_out_466;
  (* register *) pwire HA_out_467;
  (* register *) pwire HA_out_468;
  (* register *) pwire HA_out_469;
  (* register *) pwire HA_out_470;
  (* register *) pwire HA_out_471;
  (* register *) pwire HA_out_472;
  (* register *) pwire HA_out_473;
  (* register *) pwire HA_out_474;
  (* register *) pwire HA_out_475;
  (* register *) pwire HA_out_476;
  (* register *) pwire HA_out_477;
  (* register *) pwire HA_out_478;
  (* register *) pwire HA_out_479;
  (* register *) pwire HA_out_480;
  (* register *) pwire HA_out_481;
  (* register *) pwire HA_out_482;
  (* register *) pwire HA_out_483;
  (* register *) pwire HA_out_484;
  (* register *) pwire HA_out_485;
  (* register *) pwire HA_out_486;
  (* register *) pwire HA_out_487;
  (* register *) pwire HA_out_488;
  (* register *) pwire HA_out_489;
  (* register *) pwire HA_out_490;
  (* register *) pwire HA_out_491;
  (* register *) pwire HA_out_492;
  (* register *) pwire HA_out_493;
  (* register *) pwire HA_out_494;
  (* register *) pwire HA_out_495;
  (* register *) pwire HA_out_496;
  (* register *) pwire HA_out_497;
  (* register *) pwire HA_out_498;
  (* register *) pwire HA_out_499;
  (* register *) pwire HA_out_500;
  (* register *) pwire HA_out_501;
  (* register *) pwire HA_out_502;
  (* register *) pwire HA_out_503;
  (* register *) pwire HA_out_504;
  (* register *) pwire HA_out_505;
  (* register *) pwire HA_out_506;
  (* register *) pwire HA_out_507;
  (* register *) pwire HA_out_508;
  (* register *) pwire HA_out_509;
  (* register *) pwire HA_out_510;
  (* register *) pwire HA_out_511;
  (* register *) pwire HA_out_512;
  (* register *) pwire HA_out_513;
  (* register *) pwire HA_out_514;
  (* register *) pwire HA_out_515;
  (* register *) pwire HA_out_516;
  (* register *) pwire HA_out_517;
  (* register *) pwire HA_out_518;
  (* register *) pwire HA_out_519;
  (* register *) pwire HA_out_520;
  (* register *) pwire HA_out_521;
  (* register *) pwire HA_out_522;
  (* register *) pwire HA_out_523;
  (* register *) pwire HA_out_524;
  (* register *) pwire HA_out_525;
  (* register *) pwire HA_out_526;
  (* register *) pwire HA_out_527;
  (* register *) pwire HA_out_528;
  (* register *) pwire HA_out_529;
  (* register *) pwire HA_out_530;
  (* register *) pwire HA_out_531;
  (* register *) pwire HA_out_532;
  (* register *) pwire HA_out_533;
  (* register *) pwire HA_out_534;
  (* register *) pwire HA_out_535;
  (* register *) pwire HA_out_536;
  (* register *) pwire HA_out_537;
  (* register *) pwire HA_out_538;
  (* register *) pwire HA_out_539;
  (* register *) pwire HA_out_540;
  (* register *) pwire HA_out_541;
  (* register *) pwire HA_out_542;
  (* register *) pwire HA_out_543;
  (* register *) pwire HA_out_544;
  (* register *) pwire HA_out_545;
  (* register *) pwire HA_out_546;
  (* register *) pwire HA_out_547;
  (* register *) pwire HA_out_548;
  (* register *) pwire HA_out_549;
  (* register *) pwire HA_out_550;
  (* register *) pwire HA_out_551;
  (* register *) pwire HA_out_552;
  (* register *) pwire HA_out_553;
  (* register *) pwire HA_out_554;
  (* register *) pwire HA_out_555;
  (* register *) pwire HA_out_556;
  (* register *) pwire HA_out_557;
  (* register *) pwire HA_out_558;
  (* register *) pwire HA_out_559;
  (* register *) pwire HA_out_560;
  (* register *) pwire HA_out_561;
  (* register *) pwire HA_out_562;
  (* register *) pwire HA_out_563;
  (* register *) pwire HA_out_564;
  (* register *) pwire HA_out_565;
  (* register *) pwire HA_cout_0;
  (* register *) pwire HA_cout_1;
  (* register *) pwire HA_cout_2;
  (* register *) pwire HA_cout_3;
  (* register *) pwire HA_cout_4;
  (* register *) pwire HA_cout_5;
  (* register *) pwire HA_cout_6;
  (* register *) pwire HA_cout_7;
  (* register *) pwire HA_cout_8;
  (* register *) pwire HA_cout_9;
  (* register *) pwire HA_cout_10;
  (* register *) pwire HA_cout_11;
  (* register *) pwire HA_cout_12;
  (* register *) pwire HA_cout_13;
  (* register *) pwire HA_cout_14;
  (* register *) pwire HA_cout_15;
  (* register *) pwire HA_cout_16;
  (* register *) pwire HA_cout_17;
  (* register *) pwire HA_cout_18;
  (* register *) pwire HA_cout_19;
  (* register *) pwire HA_cout_20;
  (* register *) pwire HA_cout_21;
  (* register *) pwire HA_cout_22;
  (* register *) pwire HA_cout_23;
  (* register *) pwire HA_cout_24;
  (* register *) pwire HA_cout_25;
  (* register *) pwire HA_cout_26;
  (* register *) pwire HA_cout_27;
  (* register *) pwire HA_cout_28;
  (* register *) pwire HA_cout_29;
  (* register *) pwire HA_cout_30;
  (* register *) pwire HA_cout_31;
  (* register *) pwire HA_cout_32;
  (* register *) pwire HA_cout_33;
  (* register *) pwire HA_cout_34;
  (* register *) pwire HA_cout_35;
  (* register *) pwire HA_cout_36;
  (* register *) pwire HA_cout_37;
  (* register *) pwire HA_cout_38;
  (* register *) pwire HA_cout_39;
  (* register *) pwire HA_cout_40;
  (* register *) pwire HA_cout_41;
  (* register *) pwire HA_cout_42;
  (* register *) pwire HA_cout_43;
  (* register *) pwire HA_cout_44;
  (* register *) pwire HA_cout_45;
  (* register *) pwire HA_cout_46;
  (* register *) pwire HA_cout_47;
  (* register *) pwire HA_cout_48;
  (* register *) pwire HA_cout_49;
  (* register *) pwire HA_cout_50;
  (* register *) pwire HA_cout_51;
  (* register *) pwire HA_cout_52;
  (* register *) pwire HA_cout_53;
  (* register *) pwire HA_cout_54;
  (* register *) pwire HA_cout_55;
  (* register *) pwire HA_cout_56;
  (* register *) pwire HA_cout_57;
  (* register *) pwire HA_cout_58;
  (* register *) pwire HA_cout_59;
  (* register *) pwire HA_cout_60;
  (* register *) pwire HA_cout_61;
  (* register *) pwire HA_cout_62;
  (* register *) pwire HA_cout_63;
  (* register *) pwire HA_cout_64;
  (* register *) pwire HA_cout_65;
  (* register *) pwire HA_cout_66;
  (* register *) pwire HA_cout_67;
  (* register *) pwire HA_cout_68;
  (* register *) pwire HA_cout_69;
  (* register *) pwire HA_cout_70;
  (* register *) pwire HA_cout_71;
  (* register *) pwire HA_cout_72;
  (* register *) pwire HA_cout_73;
  (* register *) pwire HA_cout_74;
  (* register *) pwire HA_cout_75;
  (* register *) pwire HA_cout_76;
  (* register *) pwire HA_cout_77;
  (* register *) pwire HA_cout_78;
  (* register *) pwire HA_cout_79;
  (* register *) pwire HA_cout_80;
  (* register *) pwire HA_cout_81;
  (* register *) pwire HA_cout_82;
  (* register *) pwire HA_cout_83;
  (* register *) pwire HA_cout_84;
  (* register *) pwire HA_cout_85;
  (* register *) pwire HA_cout_86;
  (* register *) pwire HA_cout_87;
  (* register *) pwire HA_cout_88;
  (* register *) pwire HA_cout_89;
  (* register *) pwire HA_cout_90;
  (* register *) pwire HA_cout_91;
  (* register *) pwire HA_cout_92;
  (* register *) pwire HA_cout_93;
  (* register *) pwire HA_cout_94;
  (* register *) pwire HA_cout_95;
  (* register *) pwire HA_cout_96;
  (* register *) pwire HA_cout_97;
  (* register *) pwire HA_cout_98;
  (* register *) pwire HA_cout_99;
  (* register *) pwire HA_cout_100;
  (* register *) pwire HA_cout_101;
  (* register *) pwire HA_cout_102;
  (* register *) pwire HA_cout_103;
  (* register *) pwire HA_cout_104;
  (* register *) pwire HA_cout_105;
  (* register *) pwire HA_cout_106;
  (* register *) pwire HA_cout_107;
  (* register *) pwire HA_cout_108;
  (* register *) pwire HA_cout_109;
  (* register *) pwire HA_cout_110;
  (* register *) pwire HA_cout_111;
  (* register *) pwire HA_cout_112;
  (* register *) pwire HA_cout_113;
  (* register *) pwire HA_cout_114;
  (* register *) pwire HA_cout_115;
  (* register *) pwire HA_cout_116;
  (* register *) pwire HA_cout_117;
  (* register *) pwire HA_cout_118;
  (* register *) pwire HA_cout_119;
  (* register *) pwire HA_cout_120;
  (* register *) pwire HA_cout_121;
  (* register *) pwire HA_cout_122;
  (* register *) pwire HA_cout_123;
  (* register *) pwire HA_cout_124;
  (* register *) pwire HA_cout_125;
  (* register *) pwire HA_cout_126;
  (* register *) pwire HA_cout_127;
  (* register *) pwire HA_cout_128;
  (* register *) pwire HA_cout_129;
  (* register *) pwire HA_cout_130;
  (* register *) pwire HA_cout_131;
  (* register *) pwire HA_cout_132;
  (* register *) pwire HA_cout_133;
  (* register *) pwire HA_cout_134;
  (* register *) pwire HA_cout_135;
  (* register *) pwire HA_cout_136;
  (* register *) pwire HA_cout_137;
  (* register *) pwire HA_cout_138;
  (* register *) pwire HA_cout_139;
  (* register *) pwire HA_cout_140;
  (* register *) pwire HA_cout_141;
  (* register *) pwire HA_cout_142;
  (* register *) pwire HA_cout_143;
  (* register *) pwire HA_cout_144;
  (* register *) pwire HA_cout_145;
  (* register *) pwire HA_cout_146;
  (* register *) pwire HA_cout_147;
  (* register *) pwire HA_cout_148;
  (* register *) pwire HA_cout_149;
  (* register *) pwire HA_cout_150;
  (* register *) pwire HA_cout_151;
  (* register *) pwire HA_cout_152;
  (* register *) pwire HA_cout_153;
  (* register *) pwire HA_cout_154;
  (* register *) pwire HA_cout_155;
  (* register *) pwire HA_cout_156;
  (* register *) pwire HA_cout_157;
  (* register *) pwire HA_cout_158;
  (* register *) pwire HA_cout_159;
  (* register *) pwire HA_cout_160;
  (* register *) pwire HA_cout_161;
  (* register *) pwire HA_cout_162;
  (* register *) pwire HA_cout_163;
  (* register *) pwire HA_cout_164;
  (* register *) pwire HA_cout_165;
  (* register *) pwire HA_cout_166;
  (* register *) pwire HA_cout_167;
  (* register *) pwire HA_cout_168;
  (* register *) pwire HA_cout_169;
  (* register *) pwire HA_cout_170;
  (* register *) pwire HA_cout_171;
  (* register *) pwire HA_cout_172;
  (* register *) pwire HA_cout_173;
  (* register *) pwire HA_cout_174;
  (* register *) pwire HA_cout_175;
  (* register *) pwire HA_cout_176;
  (* register *) pwire HA_cout_177;
  (* register *) pwire HA_cout_178;
  (* register *) pwire HA_cout_179;
  (* register *) pwire HA_cout_180;
  (* register *) pwire HA_cout_181;
  (* register *) pwire HA_cout_182;
  (* register *) pwire HA_cout_183;
  (* register *) pwire HA_cout_184;
  (* register *) pwire HA_cout_185;
  (* register *) pwire HA_cout_186;
  (* register *) pwire HA_cout_187;
  (* register *) pwire HA_cout_188;
  (* register *) pwire HA_cout_189;
  (* register *) pwire HA_cout_190;
  (* register *) pwire HA_cout_191;
  (* register *) pwire HA_cout_192;
  (* register *) pwire HA_cout_193;
  (* register *) pwire HA_cout_194;
  (* register *) pwire HA_cout_195;
  (* register *) pwire HA_cout_196;
  (* register *) pwire HA_cout_197;
  (* register *) pwire HA_cout_198;
  (* register *) pwire HA_cout_199;
  (* register *) pwire HA_cout_200;
  (* register *) pwire HA_cout_201;
  (* register *) pwire HA_cout_202;
  (* register *) pwire HA_cout_203;
  (* register *) pwire HA_cout_204;
  (* register *) pwire HA_cout_205;
  (* register *) pwire HA_cout_206;
  (* register *) pwire HA_cout_207;
  (* register *) pwire HA_cout_208;
  (* register *) pwire HA_cout_209;
  (* register *) pwire HA_cout_210;
  (* register *) pwire HA_cout_211;
  (* register *) pwire HA_cout_212;
  (* register *) pwire HA_cout_213;
  (* register *) pwire HA_cout_214;
  (* register *) pwire HA_cout_215;
  (* register *) pwire HA_cout_216;
  (* register *) pwire HA_cout_217;
  (* register *) pwire HA_cout_218;
  (* register *) pwire HA_cout_219;
  (* register *) pwire HA_cout_220;
  (* register *) pwire HA_cout_221;
  (* register *) pwire HA_cout_222;
  (* register *) pwire HA_cout_223;
  (* register *) pwire HA_cout_224;
  (* register *) pwire HA_cout_225;
  (* register *) pwire HA_cout_226;
  (* register *) pwire HA_cout_227;
  (* register *) pwire HA_cout_228;
  (* register *) pwire HA_cout_229;
  (* register *) pwire HA_cout_230;
  (* register *) pwire HA_cout_231;
  (* register *) pwire HA_cout_232;
  (* register *) pwire HA_cout_233;
  (* register *) pwire HA_cout_234;
  (* register *) pwire HA_cout_235;
  (* register *) pwire HA_cout_236;
  (* register *) pwire HA_cout_237;
  (* register *) pwire HA_cout_238;
  (* register *) pwire HA_cout_239;
  (* register *) pwire HA_cout_240;
  (* register *) pwire HA_cout_241;
  (* register *) pwire HA_cout_242;
  (* register *) pwire HA_cout_243;
  (* register *) pwire HA_cout_244;
  (* register *) pwire HA_cout_245;
  (* register *) pwire HA_cout_246;
  (* register *) pwire HA_cout_247;
  (* register *) pwire HA_cout_248;
  (* register *) pwire HA_cout_249;
  (* register *) pwire HA_cout_250;
  (* register *) pwire HA_cout_251;
  (* register *) pwire HA_cout_252;
  (* register *) pwire HA_cout_253;
  (* register *) pwire HA_cout_254;
  (* register *) pwire HA_cout_255;
  (* register *) pwire HA_cout_256;
  (* register *) pwire HA_cout_257;
  (* register *) pwire HA_cout_258;
  (* register *) pwire HA_cout_259;
  (* register *) pwire HA_cout_260;
  (* register *) pwire HA_cout_261;
  (* register *) pwire HA_cout_262;
  (* register *) pwire HA_cout_263;
  (* register *) pwire HA_cout_264;
  (* register *) pwire HA_cout_265;
  (* register *) pwire HA_cout_266;
  (* register *) pwire HA_cout_267;
  (* register *) pwire HA_cout_268;
  (* register *) pwire HA_cout_269;
  (* register *) pwire HA_cout_270;
  (* register *) pwire HA_cout_271;
  (* register *) pwire HA_cout_272;
  (* register *) pwire HA_cout_273;
  (* register *) pwire HA_cout_274;
  (* register *) pwire HA_cout_275;
  (* register *) pwire HA_cout_276;
  (* register *) pwire HA_cout_277;
  (* register *) pwire HA_cout_278;
  (* register *) pwire HA_cout_279;
  (* register *) pwire HA_cout_280;
  (* register *) pwire HA_cout_281;
  (* register *) pwire HA_cout_282;
  (* register *) pwire HA_cout_283;
  (* register *) pwire HA_cout_284;
  (* register *) pwire HA_cout_285;
  (* register *) pwire HA_cout_286;
  (* register *) pwire HA_cout_287;
  (* register *) pwire HA_cout_288;
  (* register *) pwire HA_cout_289;
  (* register *) pwire HA_cout_290;
  (* register *) pwire HA_cout_291;
  (* register *) pwire HA_cout_292;
  (* register *) pwire HA_cout_293;
  (* register *) pwire HA_cout_294;
  (* register *) pwire HA_cout_295;
  (* register *) pwire HA_cout_296;
  (* register *) pwire HA_cout_297;
  (* register *) pwire HA_cout_298;
  (* register *) pwire HA_cout_299;
  (* register *) pwire HA_cout_300;
  (* register *) pwire HA_cout_301;
  (* register *) pwire HA_cout_302;
  (* register *) pwire HA_cout_303;
  (* register *) pwire HA_cout_304;
  (* register *) pwire HA_cout_305;
  (* register *) pwire HA_cout_306;
  (* register *) pwire HA_cout_307;
  (* register *) pwire HA_cout_308;
  (* register *) pwire HA_cout_309;
  (* register *) pwire HA_cout_310;
  (* register *) pwire HA_cout_311;
  (* register *) pwire HA_cout_312;
  (* register *) pwire HA_cout_313;
  (* register *) pwire HA_cout_314;
  (* register *) pwire HA_cout_315;
  (* register *) pwire HA_cout_316;
  (* register *) pwire HA_cout_317;
  (* register *) pwire HA_cout_318;
  (* register *) pwire HA_cout_319;
  (* register *) pwire HA_cout_320;
  (* register *) pwire HA_cout_321;
  (* register *) pwire HA_cout_322;
  (* register *) pwire HA_cout_323;
  (* register *) pwire HA_cout_324;
  (* register *) pwire HA_cout_325;
  (* register *) pwire HA_cout_326;
  (* register *) pwire HA_cout_327;
  (* register *) pwire HA_cout_328;
  (* register *) pwire HA_cout_329;
  (* register *) pwire HA_cout_330;
  (* register *) pwire HA_cout_331;
  (* register *) pwire HA_cout_332;
  (* register *) pwire HA_cout_333;
  (* register *) pwire HA_cout_334;
  (* register *) pwire HA_cout_335;
  (* register *) pwire HA_cout_336;
  (* register *) pwire HA_cout_337;
  (* register *) pwire HA_cout_338;
  (* register *) pwire HA_cout_339;
  (* register *) pwire HA_cout_340;
  (* register *) pwire HA_cout_341;
  (* register *) pwire HA_cout_342;
  (* register *) pwire HA_cout_343;
  (* register *) pwire HA_cout_344;
  (* register *) pwire HA_cout_345;
  (* register *) pwire HA_cout_346;
  (* register *) pwire HA_cout_347;
  (* register *) pwire HA_cout_348;
  (* register *) pwire HA_cout_349;
  (* register *) pwire HA_cout_350;
  (* register *) pwire HA_cout_351;
  (* register *) pwire HA_cout_352;
  (* register *) pwire HA_cout_353;
  (* register *) pwire HA_cout_354;
  (* register *) pwire HA_cout_355;
  (* register *) pwire HA_cout_356;
  (* register *) pwire HA_cout_357;
  (* register *) pwire HA_cout_358;
  (* register *) pwire HA_cout_359;
  (* register *) pwire HA_cout_360;
  (* register *) pwire HA_cout_361;
  (* register *) pwire HA_cout_362;
  (* register *) pwire HA_cout_363;
  (* register *) pwire HA_cout_364;
  (* register *) pwire HA_cout_365;
  (* register *) pwire HA_cout_366;
  (* register *) pwire HA_cout_367;
  (* register *) pwire HA_cout_368;
  (* register *) pwire HA_cout_369;
  (* register *) pwire HA_cout_370;
  (* register *) pwire HA_cout_371;
  (* register *) pwire HA_cout_372;
  (* register *) pwire HA_cout_373;
  (* register *) pwire HA_cout_374;
  (* register *) pwire HA_cout_375;
  (* register *) pwire HA_cout_376;
  (* register *) pwire HA_cout_377;
  (* register *) pwire HA_cout_378;
  (* register *) pwire HA_cout_379;
  (* register *) pwire HA_cout_380;
  (* register *) pwire HA_cout_381;
  (* register *) pwire HA_cout_382;
  (* register *) pwire HA_cout_383;
  (* register *) pwire HA_cout_384;
  (* register *) pwire HA_cout_385;
  (* register *) pwire HA_cout_386;
  (* register *) pwire HA_cout_387;
  (* register *) pwire HA_cout_388;
  (* register *) pwire HA_cout_389;
  (* register *) pwire HA_cout_390;
  (* register *) pwire HA_cout_391;
  (* register *) pwire HA_cout_392;
  (* register *) pwire HA_cout_393;
  (* register *) pwire HA_cout_394;
  (* register *) pwire HA_cout_395;
  (* register *) pwire HA_cout_396;
  (* register *) pwire HA_cout_397;
  (* register *) pwire HA_cout_398;
  (* register *) pwire HA_cout_399;
  (* register *) pwire HA_cout_400;
  (* register *) pwire HA_cout_401;
  (* register *) pwire HA_cout_402;
  (* register *) pwire HA_cout_403;
  (* register *) pwire HA_cout_404;
  (* register *) pwire HA_cout_405;
  (* register *) pwire HA_cout_406;
  (* register *) pwire HA_cout_407;
  (* register *) pwire HA_cout_408;
  (* register *) pwire HA_cout_409;
  (* register *) pwire HA_cout_410;
  (* register *) pwire HA_cout_411;
  (* register *) pwire HA_cout_412;
  (* register *) pwire HA_cout_413;
  (* register *) pwire HA_cout_414;
  (* register *) pwire HA_cout_415;
  (* register *) pwire HA_cout_416;
  (* register *) pwire HA_cout_417;
  (* register *) pwire HA_cout_418;
  (* register *) pwire HA_cout_419;
  (* register *) pwire HA_cout_420;
  (* register *) pwire HA_cout_421;
  (* register *) pwire HA_cout_422;
  (* register *) pwire HA_cout_423;
  (* register *) pwire HA_cout_424;
  (* register *) pwire HA_cout_425;
  (* register *) pwire HA_cout_426;
  (* register *) pwire HA_cout_427;
  (* register *) pwire HA_cout_428;
  (* register *) pwire HA_cout_429;
  (* register *) pwire HA_cout_430;
  (* register *) pwire HA_cout_431;
  (* register *) pwire HA_cout_432;
  (* register *) pwire HA_cout_433;
  (* register *) pwire HA_cout_434;
  (* register *) pwire HA_cout_435;
  (* register *) pwire HA_cout_436;
  (* register *) pwire HA_cout_437;
  (* register *) pwire HA_cout_438;
  (* register *) pwire HA_cout_439;
  (* register *) pwire HA_cout_440;
  (* register *) pwire HA_cout_441;
  (* register *) pwire HA_cout_442;
  (* register *) pwire HA_cout_443;
  (* register *) pwire HA_cout_444;
  (* register *) pwire HA_cout_445;
  (* register *) pwire HA_cout_446;
  (* register *) pwire HA_cout_447;
  (* register *) pwire HA_cout_448;
  (* register *) pwire HA_cout_449;
  (* register *) pwire HA_cout_450;
  (* register *) pwire HA_cout_451;
  (* register *) pwire HA_cout_452;
  (* register *) pwire HA_cout_453;
  (* register *) pwire HA_cout_454;
  (* register *) pwire HA_cout_455;
  (* register *) pwire HA_cout_456;
  (* register *) pwire HA_cout_457;
  (* register *) pwire HA_cout_458;
  (* register *) pwire HA_cout_459;
  (* register *) pwire HA_cout_460;
  (* register *) pwire HA_cout_461;
  (* register *) pwire HA_cout_462;
  (* register *) pwire HA_cout_463;
  (* register *) pwire HA_cout_464;
  (* register *) pwire HA_cout_465;
  (* register *) pwire HA_cout_466;
  (* register *) pwire HA_cout_467;
  (* register *) pwire HA_cout_468;
  (* register *) pwire HA_cout_469;
  (* register *) pwire HA_cout_470;
  (* register *) pwire HA_cout_471;
  (* register *) pwire HA_cout_472;
  (* register *) pwire HA_cout_473;
  (* register *) pwire HA_cout_474;
  (* register *) pwire HA_cout_475;
  (* register *) pwire HA_cout_476;
  (* register *) pwire HA_cout_477;
  (* register *) pwire HA_cout_478;
  (* register *) pwire HA_cout_479;
  (* register *) pwire HA_cout_480;
  (* register *) pwire HA_cout_481;
  (* register *) pwire HA_cout_482;
  (* register *) pwire HA_cout_483;
  (* register *) pwire HA_cout_484;
  (* register *) pwire HA_cout_485;
  (* register *) pwire HA_cout_486;
  (* register *) pwire HA_cout_487;
  (* register *) pwire HA_cout_488;
  (* register *) pwire HA_cout_489;
  (* register *) pwire HA_cout_490;
  (* register *) pwire HA_cout_491;
  (* register *) pwire HA_cout_492;
  (* register *) pwire HA_cout_493;
  (* register *) pwire HA_cout_494;
  (* register *) pwire HA_cout_495;
  (* register *) pwire HA_cout_496;
  (* register *) pwire HA_cout_497;
  (* register *) pwire HA_cout_498;
  (* register *) pwire HA_cout_499;
  (* register *) pwire HA_cout_500;
  (* register *) pwire HA_cout_501;
  (* register *) pwire HA_cout_502;
  (* register *) pwire HA_cout_503;
  (* register *) pwire HA_cout_504;
  (* register *) pwire HA_cout_505;
  (* register *) pwire HA_cout_506;
  (* register *) pwire HA_cout_507;
  (* register *) pwire HA_cout_508;
  (* register *) pwire HA_cout_509;
  (* register *) pwire HA_cout_510;
  (* register *) pwire HA_cout_511;
  (* register *) pwire HA_cout_512;
  (* register *) pwire HA_cout_513;
  (* register *) pwire HA_cout_514;
  (* register *) pwire HA_cout_515;
  (* register *) pwire HA_cout_516;
  (* register *) pwire HA_cout_517;
  (* register *) pwire HA_cout_518;
  (* register *) pwire HA_cout_519;
  (* register *) pwire HA_cout_520;
  (* register *) pwire HA_cout_521;
  (* register *) pwire HA_cout_522;
  (* register *) pwire HA_cout_523;
  (* register *) pwire HA_cout_524;
  (* register *) pwire HA_cout_525;
  (* register *) pwire HA_cout_526;
  (* register *) pwire HA_cout_527;
  (* register *) pwire HA_cout_528;
  (* register *) pwire HA_cout_529;
  (* register *) pwire HA_cout_530;
  (* register *) pwire HA_cout_531;
  (* register *) pwire HA_cout_532;
  (* register *) pwire HA_cout_533;
  (* register *) pwire HA_cout_534;
  (* register *) pwire HA_cout_535;
  (* register *) pwire HA_cout_536;
  (* register *) pwire HA_cout_537;
  (* register *) pwire HA_cout_538;
  (* register *) pwire HA_cout_539;
  (* register *) pwire HA_cout_540;
  (* register *) pwire HA_cout_541;
  (* register *) pwire HA_cout_542;
  (* register *) pwire HA_cout_543;
  (* register *) pwire HA_cout_544;
  (* register *) pwire HA_cout_545;
  (* register *) pwire HA_cout_546;
  (* register *) pwire HA_cout_547;
  (* register *) pwire HA_cout_548;
  (* register *) pwire HA_cout_549;
  (* register *) pwire HA_cout_550;
  (* register *) pwire HA_cout_551;
  (* register *) pwire HA_cout_552;
  (* register *) pwire HA_cout_553;
  (* register *) pwire HA_cout_554;
  (* register *) pwire HA_cout_555;
  (* register *) pwire HA_cout_556;
  (* register *) pwire HA_cout_557;
  (* register *) pwire HA_cout_558;
  (* register *) pwire HA_cout_559;
  (* register *) pwire HA_cout_560;
  (* register *) pwire HA_cout_561;
  (* register *) pwire HA_cout_562;
  (* register *) pwire HA_cout_563;
  (* register *) pwire HA_cout_564;
  (* register *) pwire HA_cout_565;
  (* register *) pwire [64:0] inp_0;

  (* register *) pwire [64:0] inp_1;

  (* register *) pwire [64:0] inp_2;

  (* register *) pwire [64:0] inp_3;

  (* register *) pwire [64:0] inp_4;

  (* register *) pwire [64:0] inp_5;

  (* register *) pwire [64:0] inp_6;

  (* register *) pwire [64:0] inp_7;

  (* register *) pwire [64:0] inp_8;

  (* register *) pwire [64:0] inp_9;

  (* register *) pwire [64:0] inp_10;

  (* register *) pwire [64:0] inp_11;

  (* register *) pwire [64:0] inp_12;

  (* register *) pwire [64:0] inp_13;

  (* register *) pwire [64:0] inp_14;

  (* register *) pwire [64:0] inp_15;

  (* register *) pwire [64:0] inp_16;

  (* register *) pwire [64:0] inp_17;

  (* register *) pwire [64:0] inp_18;

  (* register *) pwire [64:0] inp_19;

  (* register *) pwire [64:0] inp_20;

  (* register *) pwire [64:0] inp_21;

  (* register *) pwire [64:0] inp_22;

  (* register *) pwire [64:0] inp_23;

  (* register *) pwire [64:0] inp_24;

  (* register *) pwire [64:0] inp_25;

  (* register *) pwire [64:0] inp_26;

  (* register *) pwire [64:0] inp_27;

  (* register *) pwire [64:0] inp_28;

  (* register *) pwire [64:0] inp_29;

  (* register *) pwire [64:0] inp_30;

  (* register *) pwire [64:0] inp_31;

  (* register *) pwire [64:0] inp_32;

  (* register *) pwire [64:0] inp_33;

  (* register *) pwire [64:0] inp_34;

  (* register *) pwire [64:0] inp_35;

  (* register *) pwire [64:0] inp_36;

  (* register *) pwire [64:0] inp_37;

  (* register *) pwire [64:0] inp_38;

  (* register *) pwire [64:0] inp_39;

  (* register *) pwire [64:0] inp_40;

  (* register *) pwire [64:0] inp_41;

  (* register *) pwire [64:0] inp_42;

  (* register *) pwire [64:0] inp_43;

  (* register *) pwire [64:0] inp_44;

  (* register *) pwire [64:0] inp_45;

  (* register *) pwire [64:0] inp_46;

  (* register *) pwire [64:0] inp_47;

  (* register *) pwire [64:0] inp_48;

  (* register *) pwire [64:0] inp_49;

  (* register *) pwire [64:0] inp_50;

  (* register *) pwire [64:0] inp_51;

  (* register *) pwire [64:0] inp_52;

  (* register *) pwire [64:0] inp_53;

  (* register *) pwire [64:0] inp_54;

  (* register *) pwire [64:0] inp_55;

  (* register *) pwire [64:0] inp_56;

  (* register *) pwire [64:0] inp_57;

  (* register *) pwire [64:0] inp_58;

  (* register *) pwire [64:0] inp_59;

  (* register *) pwire [64:0] inp_60;

  (* register *) pwire [64:0] inp_61;

  (* register *) pwire [64:0] inp_62;

  (* register *) pwire [64:0] inp_63;

  assign inp_0[62:32]=C[62:32] & {31{R[0]}} & {31{and1}};
  assign inp_0[30:0]=C[30:0] & {31{R[0]}};
  nnXor nnXor0_31_mod(C[31],R[0],1'b1,sm_sig,inp_0[31]);
  nnXor nnXor0_63_mod(C[63],R[0],and1,sig,inp_0[63]);
  assign inp_1[62:32]=C[62:32] & {31{R[1]}} & {31{and1}};
  assign inp_1[30:0]=C[30:0] & {31{R[1]}};
  nnXor nnXor1_31_mod(C[31],R[1],1'b1,sm_sig,inp_1[31]);
  nnXor nnXor1_63_mod(C[63],R[1],and1,sig,inp_1[63]);
  assign inp_2[62:32]=C[62:32] & {31{R[2]}} & {31{and1}};
  assign inp_2[30:0]=C[30:0] & {31{R[2]}};
  nnXor nnXor2_31_mod(C[31],R[2],1'b1,sm_sig,inp_2[31]);
  nnXor nnXor2_63_mod(C[63],R[2],and1,sig,inp_2[63]);
  assign inp_3[62:32]=C[62:32] & {31{R[3]}} & {31{and1}};
  assign inp_3[30:0]=C[30:0] & {31{R[3]}};
  nnXor nnXor3_31_mod(C[31],R[3],1'b1,sm_sig,inp_3[31]);
  nnXor nnXor3_63_mod(C[63],R[3],and1,sig,inp_3[63]);
  assign inp_4[62:32]=C[62:32] & {31{R[4]}} & {31{and1}};
  assign inp_4[30:0]=C[30:0] & {31{R[4]}};
  nnXor nnXor4_31_mod(C[31],R[4],1'b1,sm_sig,inp_4[31]);
  nnXor nnXor4_63_mod(C[63],R[4],and1,sig,inp_4[63]);
  assign inp_5[62:32]=C[62:32] & {31{R[5]}} & {31{and1}};
  assign inp_5[30:0]=C[30:0] & {31{R[5]}};
  nnXor nnXor5_31_mod(C[31],R[5],1'b1,sm_sig,inp_5[31]);
  nnXor nnXor5_63_mod(C[63],R[5],and1,sig,inp_5[63]);
  assign inp_6[62:32]=C[62:32] & {31{R[6]}} & {31{and1}};
  assign inp_6[30:0]=C[30:0] & {31{R[6]}};
  nnXor nnXor6_31_mod(C[31],R[6],1'b1,sm_sig,inp_6[31]);
  nnXor nnXor6_63_mod(C[63],R[6],and1,sig,inp_6[63]);
  assign inp_7[62:32]=C[62:32] & {31{R[7]}} & {31{and1}};
  assign inp_7[30:0]=C[30:0] & {31{R[7]}};
  nnXor nnXor7_31_mod(C[31],R[7],1'b1,sm_sig,inp_7[31]);
  nnXor nnXor7_63_mod(C[63],R[7],and1,sig,inp_7[63]);
  assign inp_8[62:32]=C[62:32] & {31{R[8]}} & {31{and1}};
  assign inp_8[30:0]=C[30:0] & {31{R[8]}};
  nnXor nnXor8_31_mod(C[31],R[8],1'b1,sm_sig,inp_8[31]);
  nnXor nnXor8_63_mod(C[63],R[8],and1,sig,inp_8[63]);
  assign inp_9[62:32]=C[62:32] & {31{R[9]}} & {31{and1}};
  assign inp_9[30:0]=C[30:0] & {31{R[9]}};
  nnXor nnXor9_31_mod(C[31],R[9],1'b1,sm_sig,inp_9[31]);
  nnXor nnXor9_63_mod(C[63],R[9],and1,sig,inp_9[63]);
  assign inp_10[62:32]=C[62:32] & {31{R[10]}} & {31{and1}};
  assign inp_10[30:0]=C[30:0] & {31{R[10]}};
  nnXor nnXor10_31_mod(C[31],R[10],1'b1,sm_sig,inp_10[31]);
  nnXor nnXor10_63_mod(C[63],R[10],and1,sig,inp_10[63]);
  assign inp_11[62:32]=C[62:32] & {31{R[11]}} & {31{and1}};
  assign inp_11[30:0]=C[30:0] & {31{R[11]}};
  nnXor nnXor11_31_mod(C[31],R[11],1'b1,sm_sig,inp_11[31]);
  nnXor nnXor11_63_mod(C[63],R[11],and1,sig,inp_11[63]);
  assign inp_12[62:32]=C[62:32] & {31{R[12]}} & {31{and1}};
  assign inp_12[30:0]=C[30:0] & {31{R[12]}};
  nnXor nnXor12_31_mod(C[31],R[12],1'b1,sm_sig,inp_12[31]);
  nnXor nnXor12_63_mod(C[63],R[12],and1,sig,inp_12[63]);
  assign inp_13[62:32]=C[62:32] & {31{R[13]}} & {31{and1}};
  assign inp_13[30:0]=C[30:0] & {31{R[13]}};
  nnXor nnXor13_31_mod(C[31],R[13],1'b1,sm_sig,inp_13[31]);
  nnXor nnXor13_63_mod(C[63],R[13],and1,sig,inp_13[63]);
  assign inp_14[62:32]=C[62:32] & {31{R[14]}} & {31{and1}};
  assign inp_14[30:0]=C[30:0] & {31{R[14]}};
  nnXor nnXor14_31_mod(C[31],R[14],1'b1,sm_sig,inp_14[31]);
  nnXor nnXor14_63_mod(C[63],R[14],and1,sig,inp_14[63]);
  assign inp_15[62:32]=C[62:32] & {31{R[15]}} & {31{and1}};
  assign inp_15[30:0]=C[30:0] & {31{R[15]}};
  nnXor nnXor15_31_mod(C[31],R[15],1'b1,sm_sig,inp_15[31]);
  nnXor nnXor15_63_mod(C[63],R[15],and1,sig,inp_15[63]);
  assign inp_16[62:32]=C[62:32] & {31{R[16]}} & {31{and1}};
  assign inp_16[30:0]=C[30:0] & {31{R[16]}};
  nnXor nnXor16_31_mod(C[31],R[16],1'b1,sm_sig,inp_16[31]);
  nnXor nnXor16_63_mod(C[63],R[16],and1,sig,inp_16[63]);
  assign inp_17[62:32]=C[62:32] & {31{R[17]}} & {31{and1}};
  assign inp_17[30:0]=C[30:0] & {31{R[17]}};
  nnXor nnXor17_31_mod(C[31],R[17],1'b1,sm_sig,inp_17[31]);
  nnXor nnXor17_63_mod(C[63],R[17],and1,sig,inp_17[63]);
  assign inp_18[62:32]=C[62:32] & {31{R[18]}} & {31{and1}};
  assign inp_18[30:0]=C[30:0] & {31{R[18]}};
  nnXor nnXor18_31_mod(C[31],R[18],1'b1,sm_sig,inp_18[31]);
  nnXor nnXor18_63_mod(C[63],R[18],and1,sig,inp_18[63]);
  assign inp_19[62:32]=C[62:32] & {31{R[19]}} & {31{and1}};
  assign inp_19[30:0]=C[30:0] & {31{R[19]}};
  nnXor nnXor19_31_mod(C[31],R[19],1'b1,sm_sig,inp_19[31]);
  nnXor nnXor19_63_mod(C[63],R[19],and1,sig,inp_19[63]);
  assign inp_20[62:32]=C[62:32] & {31{R[20]}} & {31{and1}};
  assign inp_20[30:0]=C[30:0] & {31{R[20]}};
  nnXor nnXor20_31_mod(C[31],R[20],1'b1,sm_sig,inp_20[31]);
  nnXor nnXor20_63_mod(C[63],R[20],and1,sig,inp_20[63]);
  assign inp_21[62:32]=C[62:32] & {31{R[21]}} & {31{and1}};
  assign inp_21[30:0]=C[30:0] & {31{R[21]}};
  nnXor nnXor21_31_mod(C[31],R[21],1'b1,sm_sig,inp_21[31]);
  nnXor nnXor21_63_mod(C[63],R[21],and1,sig,inp_21[63]);
  assign inp_22[62:32]=C[62:32] & {31{R[22]}} & {31{and1}};
  assign inp_22[30:0]=C[30:0] & {31{R[22]}};
  nnXor nnXor22_31_mod(C[31],R[22],1'b1,sm_sig,inp_22[31]);
  nnXor nnXor22_63_mod(C[63],R[22],and1,sig,inp_22[63]);
  assign inp_23[62:32]=C[62:32] & {31{R[23]}} & {31{and1}};
  assign inp_23[30:0]=C[30:0] & {31{R[23]}};
  nnXor nnXor23_31_mod(C[31],R[23],1'b1,sm_sig,inp_23[31]);
  nnXor nnXor23_63_mod(C[63],R[23],and1,sig,inp_23[63]);
  assign inp_24[62:32]=C[62:32] & {31{R[24]}} & {31{and1}};
  assign inp_24[30:0]=C[30:0] & {31{R[24]}};
  nnXor nnXor24_31_mod(C[31],R[24],1'b1,sm_sig,inp_24[31]);
  nnXor nnXor24_63_mod(C[63],R[24],and1,sig,inp_24[63]);
  assign inp_25[62:32]=C[62:32] & {31{R[25]}} & {31{and1}};
  assign inp_25[30:0]=C[30:0] & {31{R[25]}};
  nnXor nnXor25_31_mod(C[31],R[25],1'b1,sm_sig,inp_25[31]);
  nnXor nnXor25_63_mod(C[63],R[25],and1,sig,inp_25[63]);
  assign inp_26[62:32]=C[62:32] & {31{R[26]}} & {31{and1}};
  assign inp_26[30:0]=C[30:0] & {31{R[26]}};
  nnXor nnXor26_31_mod(C[31],R[26],1'b1,sm_sig,inp_26[31]);
  nnXor nnXor26_63_mod(C[63],R[26],and1,sig,inp_26[63]);
  assign inp_27[62:32]=C[62:32] & {31{R[27]}} & {31{and1}};
  assign inp_27[30:0]=C[30:0] & {31{R[27]}};
  nnXor nnXor27_31_mod(C[31],R[27],1'b1,sm_sig,inp_27[31]);
  nnXor nnXor27_63_mod(C[63],R[27],and1,sig,inp_27[63]);
  assign inp_28[62:32]=C[62:32] & {31{R[28]}} & {31{and1}};
  assign inp_28[30:0]=C[30:0] & {31{R[28]}};
  nnXor nnXor28_31_mod(C[31],R[28],1'b1,sm_sig,inp_28[31]);
  nnXor nnXor28_63_mod(C[63],R[28],and1,sig,inp_28[63]);
  assign inp_29[62:32]=C[62:32] & {31{R[29]}} & {31{and1}};
  assign inp_29[30:0]=C[30:0] & {31{R[29]}};
  nnXor nnXor29_31_mod(C[31],R[29],1'b1,sm_sig,inp_29[31]);
  nnXor nnXor29_63_mod(C[63],R[29],and1,sig,inp_29[63]);
  assign inp_30[62:32]=C[62:32] & {31{R[30]}} & {31{and1}};
  assign inp_30[30:0]=C[30:0] & {31{R[30]}};
  nnXor nnXor30_31_mod(C[31],R[30],1'b1,sm_sig,inp_30[31]);
  nnXor nnXor30_63_mod(C[63],R[30],and1,sig,inp_30[63]);
  nnXor nnXor31_30_mod(C[30],R[31],1'b1,sm_sig,inp_31[30]);
  nnXor nnXor31_29_mod(C[29],R[31],1'b1,sm_sig,inp_31[29]);
  nnXor nnXor31_28_mod(C[28],R[31],1'b1,sm_sig,inp_31[28]);
  nnXor nnXor31_27_mod(C[27],R[31],1'b1,sm_sig,inp_31[27]);
  nnXor nnXor31_26_mod(C[26],R[31],1'b1,sm_sig,inp_31[26]);
  nnXor nnXor31_25_mod(C[25],R[31],1'b1,sm_sig,inp_31[25]);
  nnXor nnXor31_24_mod(C[24],R[31],1'b1,sm_sig,inp_31[24]);
  nnXor nnXor31_23_mod(C[23],R[31],1'b1,sm_sig,inp_31[23]);
  nnXor nnXor31_22_mod(C[22],R[31],1'b1,sm_sig,inp_31[22]);
  nnXor nnXor31_21_mod(C[21],R[31],1'b1,sm_sig,inp_31[21]);
  nnXor nnXor31_20_mod(C[20],R[31],1'b1,sm_sig,inp_31[20]);
  nnXor nnXor31_19_mod(C[19],R[31],1'b1,sm_sig,inp_31[19]);
  nnXor nnXor31_18_mod(C[18],R[31],1'b1,sm_sig,inp_31[18]);
  nnXor nnXor31_17_mod(C[17],R[31],1'b1,sm_sig,inp_31[17]);
  nnXor nnXor31_16_mod(C[16],R[31],1'b1,sm_sig,inp_31[16]);
  nnXor nnXor31_15_mod(C[15],R[31],1'b1,sm_sig,inp_31[15]);
  nnXor nnXor31_14_mod(C[14],R[31],1'b1,sm_sig,inp_31[14]);
  nnXor nnXor31_13_mod(C[13],R[31],1'b1,sm_sig,inp_31[13]);
  nnXor nnXor31_12_mod(C[12],R[31],1'b1,sm_sig,inp_31[12]);
  nnXor nnXor31_11_mod(C[11],R[31],1'b1,sm_sig,inp_31[11]);
  nnXor nnXor31_10_mod(C[10],R[31],1'b1,sm_sig,inp_31[10]);
  nnXor nnXor31_9_mod(C[9],R[31],1'b1,sm_sig,inp_31[9]);
  nnXor nnXor31_8_mod(C[8],R[31],1'b1,sm_sig,inp_31[8]);
  nnXor nnXor31_7_mod(C[7],R[31],1'b1,sm_sig,inp_31[7]);
  nnXor nnXor31_6_mod(C[6],R[31],1'b1,sm_sig,inp_31[6]);
  nnXor nnXor31_5_mod(C[5],R[31],1'b1,sm_sig,inp_31[5]);
  nnXor nnXor31_4_mod(C[4],R[31],1'b1,sm_sig,inp_31[4]);
  nnXor nnXor31_3_mod(C[3],R[31],1'b1,sm_sig,inp_31[3]);
  nnXor nnXor31_2_mod(C[2],R[31],1'b1,sm_sig,inp_31[2]);
  nnXor nnXor31_1_mod(C[1],R[31],1'b1,sm_sig,inp_31[1]);
  nnXor nnXor31_0_mod(C[0],R[31],1'b1,sm_sig,inp_31[0]);
  assign inp_31[31]=C[31] & R[31];
  assign inp_31[62:32]=C[62:32] & {31{R[31]}} &{31{and1}};
  nnXor nnXor31_63_mod(C[63],R[31],and1,sig,inp_31[63]);
  assign inp_32[62:31]=C[62:31] & {32{R[32]}} &{32{and1}};
  assign inp_32[30:0]=C[30:0] & {31{R[32]}} &{31{and1}};
  nnXor nnXor32_63_mod(C[63],R[32],and1,sig,inp_32[63]);
  assign inp_33[62:31]=C[62:31] & {32{R[33]}} &{32{and1}};
  assign inp_33[30:0]=C[30:0] & {31{R[33]}} &{31{and1}};
  nnXor nnXor33_63_mod(C[63],R[33],and1,sig,inp_33[63]);
  assign inp_34[62:31]=C[62:31] & {32{R[34]}} &{32{and1}};
  assign inp_34[30:0]=C[30:0] & {31{R[34]}} &{31{and1}};
  nnXor nnXor34_63_mod(C[63],R[34],and1,sig,inp_34[63]);
  assign inp_35[62:31]=C[62:31] & {32{R[35]}} &{32{and1}};
  assign inp_35[30:0]=C[30:0] & {31{R[35]}} &{31{and1}};
  nnXor nnXor35_63_mod(C[63],R[35],and1,sig,inp_35[63]);
  assign inp_36[62:31]=C[62:31] & {32{R[36]}} &{32{and1}};
  assign inp_36[30:0]=C[30:0] & {31{R[36]}} &{31{and1}};
  nnXor nnXor36_63_mod(C[63],R[36],and1,sig,inp_36[63]);
  assign inp_37[62:31]=C[62:31] & {32{R[37]}} &{32{and1}};
  assign inp_37[30:0]=C[30:0] & {31{R[37]}} &{31{and1}};
  nnXor nnXor37_63_mod(C[63],R[37],and1,sig,inp_37[63]);
  assign inp_38[62:31]=C[62:31] & {32{R[38]}} &{32{and1}};
  assign inp_38[30:0]=C[30:0] & {31{R[38]}} &{31{and1}};
  nnXor nnXor38_63_mod(C[63],R[38],and1,sig,inp_38[63]);
  assign inp_39[62:31]=C[62:31] & {32{R[39]}} &{32{and1}};
  assign inp_39[30:0]=C[30:0] & {31{R[39]}} &{31{and1}};
  nnXor nnXor39_63_mod(C[63],R[39],and1,sig,inp_39[63]);
  assign inp_40[62:31]=C[62:31] & {32{R[40]}} &{32{and1}};
  assign inp_40[30:0]=C[30:0] & {31{R[40]}} &{31{and1}};
  nnXor nnXor40_63_mod(C[63],R[40],and1,sig,inp_40[63]);
  assign inp_41[62:31]=C[62:31] & {32{R[41]}} &{32{and1}};
  assign inp_41[30:0]=C[30:0] & {31{R[41]}} &{31{and1}};
  nnXor nnXor41_63_mod(C[63],R[41],and1,sig,inp_41[63]);
  assign inp_42[62:31]=C[62:31] & {32{R[42]}} &{32{and1}};
  assign inp_42[30:0]=C[30:0] & {31{R[42]}} &{31{and1}};
  nnXor nnXor42_63_mod(C[63],R[42],and1,sig,inp_42[63]);
  assign inp_43[62:31]=C[62:31] & {32{R[43]}} &{32{and1}};
  assign inp_43[30:0]=C[30:0] & {31{R[43]}} &{31{and1}};
  nnXor nnXor43_63_mod(C[63],R[43],and1,sig,inp_43[63]);
  assign inp_44[62:31]=C[62:31] & {32{R[44]}} &{32{and1}};
  assign inp_44[30:0]=C[30:0] & {31{R[44]}} &{31{and1}};
  nnXor nnXor44_63_mod(C[63],R[44],and1,sig,inp_44[63]);
  assign inp_45[62:31]=C[62:31] & {32{R[45]}} &{32{and1}};
  assign inp_45[30:0]=C[30:0] & {31{R[45]}} &{31{and1}};
  nnXor nnXor45_63_mod(C[63],R[45],and1,sig,inp_45[63]);
  assign inp_46[62:31]=C[62:31] & {32{R[46]}} &{32{and1}};
  assign inp_46[30:0]=C[30:0] & {31{R[46]}} &{31{and1}};
  nnXor nnXor46_63_mod(C[63],R[46],and1,sig,inp_46[63]);
  assign inp_47[62:31]=C[62:31] & {32{R[47]}} &{32{and1}};
  assign inp_47[30:0]=C[30:0] & {31{R[47]}} &{31{and1}};
  nnXor nnXor47_63_mod(C[63],R[47],and1,sig,inp_47[63]);
  assign inp_48[62:31]=C[62:31] & {32{R[48]}} &{32{and1}};
  assign inp_48[30:0]=C[30:0] & {31{R[48]}} &{31{and1}};
  nnXor nnXor48_63_mod(C[63],R[48],and1,sig,inp_48[63]);
  assign inp_49[62:31]=C[62:31] & {32{R[49]}} &{32{and1}};
  assign inp_49[30:0]=C[30:0] & {31{R[49]}} &{31{and1}};
  nnXor nnXor49_63_mod(C[63],R[49],and1,sig,inp_49[63]);
  assign inp_50[62:31]=C[62:31] & {32{R[50]}} &{32{and1}};
  assign inp_50[30:0]=C[30:0] & {31{R[50]}} &{31{and1}};
  nnXor nnXor50_63_mod(C[63],R[50],and1,sig,inp_50[63]);
  assign inp_51[62:31]=C[62:31] & {32{R[51]}} &{32{and1}};
  assign inp_51[30:0]=C[30:0] & {31{R[51]}} &{31{and1}};
  nnXor nnXor51_63_mod(C[63],R[51],and1,sig,inp_51[63]);
  assign inp_52[62:31]=C[62:31] & {32{R[52]}} &{32{and1}};
  assign inp_52[30:0]=C[30:0] & {31{R[52]}} &{31{and1}};
  nnXor nnXor52_63_mod(C[63],R[52],and1,sig,inp_52[63]);
  assign inp_53[62:31]=C[62:31] & {32{R[53]}} &{32{and1}};
  assign inp_53[30:0]=C[30:0] & {31{R[53]}} &{31{and1}};
  nnXor nnXor53_63_mod(C[63],R[53],and1,sig,inp_53[63]);
  assign inp_54[62:31]=C[62:31] & {32{R[54]}} &{32{and1}};
  assign inp_54[30:0]=C[30:0] & {31{R[54]}} &{31{and1}};
  nnXor nnXor54_63_mod(C[63],R[54],and1,sig,inp_54[63]);
  assign inp_55[62:31]=C[62:31] & {32{R[55]}} &{32{and1}};
  assign inp_55[30:0]=C[30:0] & {31{R[55]}} &{31{and1}};
  nnXor nnXor55_63_mod(C[63],R[55],and1,sig,inp_55[63]);
  assign inp_56[62:31]=C[62:31] & {32{R[56]}} &{32{and1}};
  assign inp_56[30:0]=C[30:0] & {31{R[56]}} &{31{and1}};
  nnXor nnXor56_63_mod(C[63],R[56],and1,sig,inp_56[63]);
  assign inp_57[62:31]=C[62:31] & {32{R[57]}} &{32{and1}};
  assign inp_57[30:0]=C[30:0] & {31{R[57]}} &{31{and1}};
  nnXor nnXor57_63_mod(C[63],R[57],and1,sig,inp_57[63]);
  assign inp_58[62:31]=C[62:31] & {32{R[58]}} &{32{and1}};
  assign inp_58[30:0]=C[30:0] & {31{R[58]}} &{31{and1}};
  nnXor nnXor58_63_mod(C[63],R[58],and1,sig,inp_58[63]);
  assign inp_59[62:31]=C[62:31] & {32{R[59]}} &{32{and1}};
  assign inp_59[30:0]=C[30:0] & {31{R[59]}} &{31{and1}};
  nnXor nnXor59_63_mod(C[63],R[59],and1,sig,inp_59[63]);
  assign inp_60[62:31]=C[62:31] & {32{R[60]}} &{32{and1}};
  assign inp_60[30:0]=C[30:0] & {31{R[60]}} &{31{and1}};
  nnXor nnXor60_63_mod(C[63],R[60],and1,sig,inp_60[63]);
  assign inp_61[62:31]=C[62:31] & {32{R[61]}} &{32{and1}};
  assign inp_61[30:0]=C[30:0] & {31{R[61]}} &{31{and1}};
  nnXor nnXor61_63_mod(C[63],R[61],and1,sig,inp_61[63]);
  assign inp_62[62:31]=C[62:31] & {32{R[62]}} &{32{and1}};
  assign inp_62[30:0]=C[30:0] & {31{R[62]}} &{31{and1}};
  nnXor nnXor62_63_mod(C[63],R[62],and1,sig,inp_62[63]);
  assign inp_63[63]=C[63] & R[63] & and1;
  nnXor nnXor63_62_mod(C[62],R[63],and1,sig,inp_63[62]);
  nnXor nnXor63_61_mod(C[61],R[63],and1,sig,inp_63[61]);
  nnXor nnXor63_60_mod(C[60],R[63],and1,sig,inp_63[60]);
  nnXor nnXor63_59_mod(C[59],R[63],and1,sig,inp_63[59]);
  nnXor nnXor63_58_mod(C[58],R[63],and1,sig,inp_63[58]);
  nnXor nnXor63_57_mod(C[57],R[63],and1,sig,inp_63[57]);
  nnXor nnXor63_56_mod(C[56],R[63],and1,sig,inp_63[56]);
  nnXor nnXor63_55_mod(C[55],R[63],and1,sig,inp_63[55]);
  nnXor nnXor63_54_mod(C[54],R[63],and1,sig,inp_63[54]);
  nnXor nnXor63_53_mod(C[53],R[63],and1,sig,inp_63[53]);
  nnXor nnXor63_52_mod(C[52],R[63],and1,sig,inp_63[52]);
  nnXor nnXor63_51_mod(C[51],R[63],and1,sig,inp_63[51]);
  nnXor nnXor63_50_mod(C[50],R[63],and1,sig,inp_63[50]);
  nnXor nnXor63_49_mod(C[49],R[63],and1,sig,inp_63[49]);
  nnXor nnXor63_48_mod(C[48],R[63],and1,sig,inp_63[48]);
  nnXor nnXor63_47_mod(C[47],R[63],and1,sig,inp_63[47]);
  nnXor nnXor63_46_mod(C[46],R[63],and1,sig,inp_63[46]);
  nnXor nnXor63_45_mod(C[45],R[63],and1,sig,inp_63[45]);
  nnXor nnXor63_44_mod(C[44],R[63],and1,sig,inp_63[44]);
  nnXor nnXor63_43_mod(C[43],R[63],and1,sig,inp_63[43]);
  nnXor nnXor63_42_mod(C[42],R[63],and1,sig,inp_63[42]);
  nnXor nnXor63_41_mod(C[41],R[63],and1,sig,inp_63[41]);
  nnXor nnXor63_40_mod(C[40],R[63],and1,sig,inp_63[40]);
  nnXor nnXor63_39_mod(C[39],R[63],and1,sig,inp_63[39]);
  nnXor nnXor63_38_mod(C[38],R[63],and1,sig,inp_63[38]);
  nnXor nnXor63_37_mod(C[37],R[63],and1,sig,inp_63[37]);
  nnXor nnXor63_36_mod(C[36],R[63],and1,sig,inp_63[36]);
  nnXor nnXor63_35_mod(C[35],R[63],and1,sig,inp_63[35]);
  nnXor nnXor63_34_mod(C[34],R[63],and1,sig,inp_63[34]);
  nnXor nnXor63_33_mod(C[33],R[63],and1,sig,inp_63[33]);
  nnXor nnXor63_32_mod(C[32],R[63],and1,sig,inp_63[32]);
  nnXor nnXor63_31_mod(C[31],R[63],and1,sig,inp_63[31]);
  nnXor nnXor63_30_mod(C[30],R[63],and1,sig,inp_63[30]);
  nnXor nnXor63_29_mod(C[29],R[63],and1,sig,inp_63[29]);
  nnXor nnXor63_28_mod(C[28],R[63],and1,sig,inp_63[28]);
  nnXor nnXor63_27_mod(C[27],R[63],and1,sig,inp_63[27]);
  nnXor nnXor63_26_mod(C[26],R[63],and1,sig,inp_63[26]);
  nnXor nnXor63_25_mod(C[25],R[63],and1,sig,inp_63[25]);
  nnXor nnXor63_24_mod(C[24],R[63],and1,sig,inp_63[24]);
  nnXor nnXor63_23_mod(C[23],R[63],and1,sig,inp_63[23]);
  nnXor nnXor63_22_mod(C[22],R[63],and1,sig,inp_63[22]);
  nnXor nnXor63_21_mod(C[21],R[63],and1,sig,inp_63[21]);
  nnXor nnXor63_20_mod(C[20],R[63],and1,sig,inp_63[20]);
  nnXor nnXor63_19_mod(C[19],R[63],and1,sig,inp_63[19]);
  nnXor nnXor63_18_mod(C[18],R[63],and1,sig,inp_63[18]);
  nnXor nnXor63_17_mod(C[17],R[63],and1,sig,inp_63[17]);
  nnXor nnXor63_16_mod(C[16],R[63],and1,sig,inp_63[16]);
  nnXor nnXor63_15_mod(C[15],R[63],and1,sig,inp_63[15]);
  nnXor nnXor63_14_mod(C[14],R[63],and1,sig,inp_63[14]);
  nnXor nnXor63_13_mod(C[13],R[63],and1,sig,inp_63[13]);
  nnXor nnXor63_12_mod(C[12],R[63],and1,sig,inp_63[12]);
  nnXor nnXor63_11_mod(C[11],R[63],and1,sig,inp_63[11]);
  nnXor nnXor63_10_mod(C[10],R[63],and1,sig,inp_63[10]);
  nnXor nnXor63_9_mod(C[9],R[63],and1,sig,inp_63[9]);
  nnXor nnXor63_8_mod(C[8],R[63],and1,sig,inp_63[8]);
  nnXor nnXor63_7_mod(C[7],R[63],and1,sig,inp_63[7]);
  nnXor nnXor63_6_mod(C[6],R[63],and1,sig,inp_63[6]);
  nnXor nnXor63_5_mod(C[5],R[63],and1,sig,inp_63[5]);
  nnXor nnXor63_4_mod(C[4],R[63],and1,sig,inp_63[4]);
  nnXor nnXor63_3_mod(C[3],R[63],and1,sig,inp_63[3]);
  nnXor nnXor63_2_mod(C[2],R[63],and1,sig,inp_63[2]);
  nnXor nnXor63_1_mod(C[1],R[63],and1,sig,inp_63[1]);
  nnXor nnXor63_0_mod(C[0],R[63],and1,sig,inp_63[0]);
  assign A_out[0]=REGS_1893;
  assign A_out[1]=REGS_1894;
  assign A_out[2]=REGS_1895;
  assign A_out[3]=REGS_1896;
  assign A_out[4]=REGS_1897;
  assign A_out[5]=REGS_1898;
  assign A_out[6]=REGS_1899;
  assign A_out[7]=HA_out_267;
  assign A_out[8]=HA_out_315;
  assign A_out[9]=HA_out_369;
  assign A_out[10]=HA_out_447;
  assign A_out[11]=HA_cout_447;
  assign A_out[12]=HA_cout_448;
  assign A_out[13]=HA_cout_449;
  assign A_out[14]=HA_cout_450;
  assign A_out[15]=HA_cout_451;
  assign A_out[16]=HA_cout_452;
  assign A_out[17]=HA_cout_453;
  assign A_out[18]=HA_cout_454;
  assign A_out[19]=HA_cout_455;
  assign A_out[20]=HA_cout_456;
  assign A_out[21]=HA_cout_457;
  assign A_out[22]=HA_cout_458;
  assign A_out[23]=HA_cout_459;
  assign A_out[24]=HA_cout_460;
  assign A_out[25]=HA_cout_461;
  assign A_out[26]=HA_cout_462;
  assign A_out[27]=HA_cout_463;
  assign A_out[28]=HA_cout_464;
  assign A_out[29]=HA_cout_465;
  assign A_out[30]=HA_cout_466;
  assign A_out[31]=HA_cout_467;
  assign A_out[32]=HA_cout_468;
  assign A_out[33]=HA_cout_469;
  assign A_out[34]=HA_cout_470;
  assign A_out[35]=HA_cout_471;
  assign A_out[36]=HA_cout_472;
  assign A_out[37]=HA_cout_473;
  assign A_out[38]=HA_cout_474;
  assign A_out[39]=HA_cout_475;
  assign A_out[40]=HA_cout_476;
  assign A_out[41]=HA_cout_477;
  assign A_out[42]=HA_cout_478;
  assign A_out[43]=HA_cout_479;
  assign A_out[44]=HA_cout_480;
  assign A_out[45]=HA_cout_481;
  assign A_out[46]=HA_cout_482;
  assign A_out[47]=HA_cout_483;
  assign A_out[48]=HA_cout_484;
  assign A_out[49]=HA_cout_485;
  assign A_out[50]=HA_cout_486;
  assign A_out[51]=HA_cout_487;
  assign A_out[52]=HA_cout_488;
  assign A_out[53]=HA_cout_489;
  assign A_out[54]=HA_cout_490;
  assign A_out[55]=HA_cout_491;
  assign A_out[56]=HA_cout_492;
  assign A_out[57]=HA_cout_493;
  assign A_out[58]=HA_cout_494;
  assign A_out[59]=HA_cout_495;
  assign A_out[60]=HA_cout_496;
  assign A_out[61]=HA_cout_497;
  assign A_out[62]=HA_cout_498;
  assign A_out[63]=HA_cout_499;
  assign A_out[64]=HA_cout_500;
  assign A_out[65]=HA_cout_501;
  assign A_out[66]=HA_cout_502;
  assign A_out[67]=HA_cout_503;
  assign A_out[68]=FA_cout_3844;
  assign A_out[69]=FA_cout_3845;
  assign A_out[70]=HA_cout_504;
  assign A_out[71]=HA_cout_505;
  assign A_out[72]=HA_cout_506;
  assign A_out[73]=HA_cout_507;
  assign A_out[74]=HA_cout_508;
  assign B_out[11]=HA_out_448;
  assign B_out[12]=HA_out_449;
  assign B_out[13]=HA_out_450;
  assign B_out[14]=HA_out_451;
  assign B_out[15]=HA_out_452;
  assign B_out[16]=HA_out_453;
  assign B_out[17]=HA_out_454;
  assign B_out[18]=HA_out_455;
  assign B_out[19]=HA_out_456;
  assign B_out[20]=HA_out_457;
  assign B_out[21]=HA_out_458;
  assign B_out[22]=HA_out_459;
  assign B_out[23]=HA_out_460;
  assign B_out[24]=HA_out_461;
  assign B_out[25]=HA_out_462;
  assign B_out[26]=HA_out_463;
  assign B_out[27]=HA_out_464;
  assign B_out[28]=HA_out_465;
  assign B_out[29]=HA_out_466;
  assign B_out[30]=HA_out_467;
  assign B_out[31]=HA_out_468;
  assign B_out[32]=HA_out_469;
  assign B_out[33]=HA_out_470;
  assign B_out[34]=HA_out_471;
  assign B_out[35]=HA_out_472;
  assign B_out[36]=HA_out_473;
  assign B_out[37]=HA_out_474;
  assign B_out[38]=HA_out_475;
  assign B_out[39]=HA_out_476;
  assign B_out[40]=HA_out_477;
  assign B_out[41]=HA_out_478;
  assign B_out[42]=HA_out_479;
  assign B_out[43]=HA_out_480;
  assign B_out[44]=HA_out_481;
  assign B_out[45]=HA_out_482;
  assign B_out[46]=HA_out_483;
  assign B_out[47]=HA_out_484;
  assign B_out[48]=HA_out_485;
  assign B_out[49]=HA_out_486;
  assign B_out[50]=HA_out_487;
  assign B_out[51]=HA_out_488;
  assign B_out[52]=HA_out_489;
  assign B_out[53]=HA_out_490;
  assign B_out[54]=HA_out_491;
  assign B_out[55]=HA_out_492;
  assign B_out[56]=HA_out_493;
  assign B_out[57]=HA_out_494;
  assign B_out[58]=HA_out_495;
  assign B_out[59]=HA_out_496;
  assign B_out[60]=HA_out_497;
  assign B_out[61]=HA_out_498;
  assign B_out[62]=HA_out_499;
  assign B_out[63]=HA_out_500;
  assign B_out[64]=HA_out_501;
  assign B_out[65]=HA_out_502;
  assign B_out[66]=HA_out_503;
  assign B_out[67]=FA_out_3844;
  assign B_out[68]=FA_out_3845;
  assign B_out[69]=HA_out_504;
  assign B_out[70]=HA_out_505;
  assign B_out[71]=HA_out_506;
  assign B_out[72]=HA_out_507;
  assign B_out[73]=HA_out_508;
  assign B_out[74]=HA_out_509;
  assign A_out[75]=HA_cout_509;
  assign B_out[75]=HA_out_510;
  assign A_out[76]=HA_cout_510;
  assign B_out[76]=HA_out_511;
  assign A_out[77]=HA_cout_511;
  assign B_out[77]=HA_out_512;
  assign A_out[78]=HA_cout_512;
  assign B_out[78]=HA_out_513;
  assign A_out[79]=HA_cout_513;
  assign B_out[79]=HA_out_514;
  assign A_out[80]=HA_cout_514;
  assign B_out[80]=HA_out_515;
  assign A_out[81]=HA_cout_515;
  assign B_out[81]=HA_out_516;
  assign A_out[82]=HA_cout_516;
  assign B_out[82]=HA_out_517;
  assign A_out[83]=HA_cout_517;
  assign B_out[83]=HA_out_518;
  assign A_out[84]=HA_cout_518;
  assign B_out[84]=HA_out_519;
  assign A_out[85]=HA_cout_519;
  assign B_out[85]=HA_out_520;
  assign A_out[86]=HA_cout_520;
  assign B_out[86]=HA_out_521;
  assign A_out[87]=HA_cout_521;
  assign B_out[87]=HA_out_522;
  assign A_out[88]=HA_cout_522;
  assign B_out[88]=HA_out_523;
  assign A_out[89]=HA_cout_523;
  assign B_out[89]=HA_out_524;
  assign A_out[90]=HA_cout_524;
  assign B_out[90]=HA_out_525;
  assign A_out[91]=HA_cout_525;
  assign B_out[91]=HA_out_526;
  assign A_out[92]=HA_cout_526;
  assign B_out[92]=HA_out_527;
  assign A_out[93]=HA_cout_527;
  assign B_out[93]=HA_out_528;
  assign A_out[94]=HA_cout_528;
  assign B_out[94]=HA_out_529;
  assign A_out[95]=HA_cout_529;
  assign B_out[95]=HA_out_530;
  assign A_out[96]=HA_cout_530;
  assign B_out[96]=HA_out_531;
  assign A_out[97]=HA_cout_531;
  assign B_out[97]=HA_out_532;
  assign A_out[98]=HA_cout_532;
  assign B_out[98]=HA_out_533;
  assign A_out[99]=HA_cout_533;
  assign B_out[99]=HA_out_534;
  assign A_out[100]=HA_cout_534;
  assign B_out[100]=HA_out_535;
  assign A_out[101]=HA_cout_535;
  assign B_out[101]=HA_out_536;
  assign A_out[102]=HA_cout_536;
  assign B_out[102]=HA_out_537;
  assign A_out[103]=HA_cout_537;
  assign B_out[103]=HA_out_538;
  assign A_out[104]=HA_cout_538;
  assign B_out[104]=HA_out_539;
  assign A_out[105]=HA_cout_539;
  assign B_out[105]=HA_out_540;
  assign A_out[106]=HA_cout_540;
  assign B_out[106]=HA_out_541;
  assign A_out[107]=HA_cout_541;
  assign B_out[107]=HA_out_542;
  assign A_out[108]=HA_cout_542;
  assign B_out[108]=HA_out_543;
  assign A_out[109]=HA_cout_543;
  assign B_out[109]=HA_out_544;
  assign A_out[110]=HA_cout_544;
  assign B_out[110]=HA_out_545;
  assign A_out[111]=HA_cout_545;
  assign B_out[111]=HA_out_546;
  assign A_out[112]=HA_cout_546;
  assign B_out[112]=HA_out_547;
  assign A_out[113]=HA_cout_547;
  assign B_out[113]=HA_out_548;
  assign A_out[114]=HA_cout_548;
  assign B_out[114]=HA_out_549;
  assign A_out[115]=HA_cout_549;
  assign B_out[115]=HA_out_550;
  assign A_out[116]=HA_cout_550;
  assign B_out[116]=HA_out_551;
  assign A_out[117]=HA_cout_551;
  assign B_out[117]=HA_out_552;
  assign A_out[118]=HA_cout_552;
  assign B_out[118]=HA_out_553;
  assign A_out[119]=HA_cout_553;
  assign B_out[119]=HA_out_554;
  assign A_out[120]=HA_cout_554;
  assign B_out[120]=HA_out_555;
  assign A_out[121]=HA_cout_555;
  assign B_out[121]=HA_out_556;
  assign A_out[122]=HA_cout_556;
  assign B_out[122]=HA_out_557;
  assign A_out[123]=HA_cout_557;
  assign B_out[123]=HA_out_558;
  assign A_out[124]=HA_cout_558;
  assign B_out[124]=HA_out_559;
  assign A_out[125]=HA_cout_559;
  assign B_out[125]=HA_out_560;
  assign A_out[126]=HA_cout_560;
  assign B_out[126]=HA_out_561;
  assign A_out[127]=HA_cout_561;
  assign B_out[127]=HA_out_562;
  assign B_out[0]=1'b0;
  assign B_out[1]=1'b0;
  assign B_out[2]=1'b0;
  assign B_out[3]=1'b0;
  assign B_out[4]=1'b0;
  assign B_out[5]=1'b0;
  assign B_out[6]=1'b0;
  assign B_out[7]=1'b0;
  assign B_out[8]=1'b0;
  assign B_out[9]=1'b0;
  assign B_out[10]=1'b0;

  assign {FA_cout_0,FA_out_0}=inp_0[2]+inp_1[1]+inp_2[0];
  assign {FA_cout_1,FA_out_1}=inp_0[3]+inp_1[2]+inp_2[1];
  assign {FA_cout_2,FA_out_2}=inp_0[4]+inp_1[3]+inp_2[2];
  assign {FA_cout_3,FA_out_3}=inp_0[5]+inp_1[4]+inp_2[3];
  assign {FA_cout_4,FA_out_4}=inp_0[6]+inp_1[5]+inp_2[4];
  assign {FA_cout_5,FA_out_5}=inp_0[7]+inp_1[6]+inp_2[5];
  assign {FA_cout_6,FA_out_6}=inp_0[8]+inp_1[7]+inp_2[6];
  assign {FA_cout_7,FA_out_7}=inp_0[9]+inp_1[8]+inp_2[7];
  assign {FA_cout_8,FA_out_8}=inp_0[10]+inp_1[9]+inp_2[8];
  assign {FA_cout_9,FA_out_9}=inp_0[11]+inp_1[10]+inp_2[9];
  assign {FA_cout_10,FA_out_10}=inp_0[12]+inp_1[11]+inp_2[10];
  assign {FA_cout_11,FA_out_11}=inp_0[13]+inp_1[12]+inp_2[11];
  assign {FA_cout_12,FA_out_12}=inp_0[14]+inp_1[13]+inp_2[12];
  assign {FA_cout_13,FA_out_13}=inp_0[15]+inp_1[14]+inp_2[13];
  assign {FA_cout_14,FA_out_14}=inp_0[16]+inp_1[15]+inp_2[14];
  assign {FA_cout_15,FA_out_15}=inp_0[17]+inp_1[16]+inp_2[15];
  assign {FA_cout_16,FA_out_16}=inp_0[18]+inp_1[17]+inp_2[16];
  assign {FA_cout_17,FA_out_17}=inp_0[19]+inp_1[18]+inp_2[17];
  assign {FA_cout_18,FA_out_18}=inp_0[20]+inp_1[19]+inp_2[18];
  assign {FA_cout_19,FA_out_19}=inp_0[21]+inp_1[20]+inp_2[19];
  assign {FA_cout_20,FA_out_20}=inp_0[22]+inp_1[21]+inp_2[20];
  assign {FA_cout_21,FA_out_21}=inp_0[23]+inp_1[22]+inp_2[21];
  assign {FA_cout_22,FA_out_22}=inp_0[24]+inp_1[23]+inp_2[22];
  assign {FA_cout_23,FA_out_23}=inp_0[25]+inp_1[24]+inp_2[23];
  assign {FA_cout_24,FA_out_24}=inp_0[26]+inp_1[25]+inp_2[24];
  assign {FA_cout_25,FA_out_25}=inp_0[27]+inp_1[26]+inp_2[25];
  assign {FA_cout_26,FA_out_26}=inp_0[28]+inp_1[27]+inp_2[26];
  assign {FA_cout_27,FA_out_27}=inp_0[29]+inp_1[28]+inp_2[27];
  assign {FA_cout_28,FA_out_28}=inp_0[30]+inp_1[29]+inp_2[28];
  assign {FA_cout_29,FA_out_29}=inp_0[31]+inp_1[30]+inp_2[29];
  assign {FA_cout_30,FA_out_30}=inp_0[32]+inp_1[31]+inp_2[30];
  assign {FA_cout_31,FA_out_31}=inp_0[33]+inp_1[32]+inp_2[31];
  assign {FA_cout_32,FA_out_32}=inp_0[34]+inp_1[33]+inp_2[32];
  assign {FA_cout_33,FA_out_33}=inp_0[35]+inp_1[34]+inp_2[33];
  assign {FA_cout_34,FA_out_34}=inp_0[36]+inp_1[35]+inp_2[34];
  assign {FA_cout_35,FA_out_35}=inp_0[37]+inp_1[36]+inp_2[35];
  assign {FA_cout_36,FA_out_36}=inp_0[38]+inp_1[37]+inp_2[36];
  assign {FA_cout_37,FA_out_37}=inp_0[39]+inp_1[38]+inp_2[37];
  assign {FA_cout_38,FA_out_38}=inp_0[40]+inp_1[39]+inp_2[38];
  assign {FA_cout_39,FA_out_39}=inp_0[41]+inp_1[40]+inp_2[39];
  assign {FA_cout_40,FA_out_40}=inp_0[42]+inp_1[41]+inp_2[40];
  assign {FA_cout_41,FA_out_41}=inp_0[43]+inp_1[42]+inp_2[41];
  assign {FA_cout_42,FA_out_42}=inp_0[44]+inp_1[43]+inp_2[42];
  assign {FA_cout_43,FA_out_43}=inp_0[45]+inp_1[44]+inp_2[43];
  assign {FA_cout_44,FA_out_44}=inp_0[46]+inp_1[45]+inp_2[44];
  assign {FA_cout_45,FA_out_45}=inp_0[47]+inp_1[46]+inp_2[45];
  assign {FA_cout_46,FA_out_46}=inp_0[48]+inp_1[47]+inp_2[46];
  assign {FA_cout_47,FA_out_47}=inp_0[49]+inp_1[48]+inp_2[47];
  assign {FA_cout_48,FA_out_48}=inp_0[50]+inp_1[49]+inp_2[48];
  assign {FA_cout_49,FA_out_49}=inp_0[51]+inp_1[50]+inp_2[49];
  assign {FA_cout_50,FA_out_50}=inp_0[52]+inp_1[51]+inp_2[50];
  assign {FA_cout_51,FA_out_51}=inp_0[53]+inp_1[52]+inp_2[51];
  assign {FA_cout_52,FA_out_52}=inp_0[54]+inp_1[53]+inp_2[52];
  assign {FA_cout_53,FA_out_53}=inp_0[55]+inp_1[54]+inp_2[53];
  assign {FA_cout_54,FA_out_54}=inp_0[56]+inp_1[55]+inp_2[54];
  assign {FA_cout_55,FA_out_55}=inp_0[57]+inp_1[56]+inp_2[55];
  assign {FA_cout_56,FA_out_56}=inp_0[58]+inp_1[57]+inp_2[56];
  assign {FA_cout_57,FA_out_57}=inp_0[59]+inp_1[58]+inp_2[57];
  assign {FA_cout_58,FA_out_58}=inp_0[60]+inp_1[59]+inp_2[58];
  assign {FA_cout_59,FA_out_59}=inp_0[61]+inp_1[60]+inp_2[59];
  assign {FA_cout_60,FA_out_60}=inp_0[62]+inp_1[61]+inp_2[60];
  assign {FA_cout_61,FA_out_61}=inp_0[63]+inp_1[62]+inp_2[61];
  assign {FA_cout_62,FA_out_62}=sig+inp_1[63]+inp_2[62];
  assign {FA_cout_63,FA_out_63}=inp_2[63]+inp_3[62]+inp_4[61];
  assign {FA_cout_64,FA_out_64}=inp_3[2]+inp_4[1]+inp_5[0];
  assign {FA_cout_65,FA_out_65}=inp_3[3]+inp_4[2]+inp_5[1];
  assign {FA_cout_66,FA_out_66}=inp_3[4]+inp_4[3]+inp_5[2];
  assign {FA_cout_67,FA_out_67}=inp_3[5]+inp_4[4]+inp_5[3];
  assign {FA_cout_68,FA_out_68}=inp_3[6]+inp_4[5]+inp_5[4];
  assign {FA_cout_69,FA_out_69}=inp_3[7]+inp_4[6]+inp_5[5];
  assign {FA_cout_70,FA_out_70}=inp_3[8]+inp_4[7]+inp_5[6];
  assign {FA_cout_71,FA_out_71}=inp_3[9]+inp_4[8]+inp_5[7];
  assign {FA_cout_72,FA_out_72}=inp_3[10]+inp_4[9]+inp_5[8];
  assign {FA_cout_73,FA_out_73}=inp_3[11]+inp_4[10]+inp_5[9];
  assign {FA_cout_74,FA_out_74}=inp_3[12]+inp_4[11]+inp_5[10];
  assign {FA_cout_75,FA_out_75}=inp_3[13]+inp_4[12]+inp_5[11];
  assign {FA_cout_76,FA_out_76}=inp_3[14]+inp_4[13]+inp_5[12];
  assign {FA_cout_77,FA_out_77}=inp_3[15]+inp_4[14]+inp_5[13];
  assign {FA_cout_78,FA_out_78}=inp_3[16]+inp_4[15]+inp_5[14];
  assign {FA_cout_79,FA_out_79}=inp_3[17]+inp_4[16]+inp_5[15];
  assign {FA_cout_80,FA_out_80}=inp_3[18]+inp_4[17]+inp_5[16];
  assign {FA_cout_81,FA_out_81}=inp_3[19]+inp_4[18]+inp_5[17];
  assign {FA_cout_82,FA_out_82}=inp_3[20]+inp_4[19]+inp_5[18];
  assign {FA_cout_83,FA_out_83}=inp_3[21]+inp_4[20]+inp_5[19];
  assign {FA_cout_84,FA_out_84}=inp_3[22]+inp_4[21]+inp_5[20];
  assign {FA_cout_85,FA_out_85}=inp_3[23]+inp_4[22]+inp_5[21];
  assign {FA_cout_86,FA_out_86}=inp_3[24]+inp_4[23]+inp_5[22];
  assign {FA_cout_87,FA_out_87}=inp_3[25]+inp_4[24]+inp_5[23];
  assign {FA_cout_88,FA_out_88}=inp_3[26]+inp_4[25]+inp_5[24];
  assign {FA_cout_89,FA_out_89}=inp_3[27]+inp_4[26]+inp_5[25];
  assign {FA_cout_90,FA_out_90}=inp_3[28]+inp_4[27]+inp_5[26];
  assign {FA_cout_91,FA_out_91}=inp_3[29]+inp_4[28]+inp_5[27];
  assign {FA_cout_92,FA_out_92}=inp_3[30]+inp_4[29]+inp_5[28];
  assign {FA_cout_93,FA_out_93}=inp_3[31]+inp_4[30]+inp_5[29];
  assign {FA_cout_94,FA_out_94}=inp_3[32]+inp_4[31]+inp_5[30];
  assign {FA_cout_95,FA_out_95}=inp_3[33]+inp_4[32]+inp_5[31];
  assign {FA_cout_96,FA_out_96}=inp_3[34]+inp_4[33]+inp_5[32];
  assign {FA_cout_97,FA_out_97}=inp_3[35]+inp_4[34]+inp_5[33];
  assign {FA_cout_98,FA_out_98}=inp_3[36]+inp_4[35]+inp_5[34];
  assign {FA_cout_99,FA_out_99}=inp_3[37]+inp_4[36]+inp_5[35];
  assign {FA_cout_100,FA_out_100}=inp_3[38]+inp_4[37]+inp_5[36];
  assign {FA_cout_101,FA_out_101}=inp_3[39]+inp_4[38]+inp_5[37];
  assign {FA_cout_102,FA_out_102}=inp_3[40]+inp_4[39]+inp_5[38];
  assign {FA_cout_103,FA_out_103}=inp_3[41]+inp_4[40]+inp_5[39];
  assign {FA_cout_104,FA_out_104}=inp_3[42]+inp_4[41]+inp_5[40];
  assign {FA_cout_105,FA_out_105}=inp_3[43]+inp_4[42]+inp_5[41];
  assign {FA_cout_106,FA_out_106}=inp_3[44]+inp_4[43]+inp_5[42];
  assign {FA_cout_107,FA_out_107}=inp_3[45]+inp_4[44]+inp_5[43];
  assign {FA_cout_108,FA_out_108}=inp_3[46]+inp_4[45]+inp_5[44];
  assign {FA_cout_109,FA_out_109}=inp_3[47]+inp_4[46]+inp_5[45];
  assign {FA_cout_110,FA_out_110}=inp_3[48]+inp_4[47]+inp_5[46];
  assign {FA_cout_111,FA_out_111}=inp_3[49]+inp_4[48]+inp_5[47];
  assign {FA_cout_112,FA_out_112}=inp_3[50]+inp_4[49]+inp_5[48];
  assign {FA_cout_113,FA_out_113}=inp_3[51]+inp_4[50]+inp_5[49];
  assign {FA_cout_114,FA_out_114}=inp_3[52]+inp_4[51]+inp_5[50];
  assign {FA_cout_115,FA_out_115}=inp_3[53]+inp_4[52]+inp_5[51];
  assign {FA_cout_116,FA_out_116}=inp_3[54]+inp_4[53]+inp_5[52];
  assign {FA_cout_117,FA_out_117}=inp_3[55]+inp_4[54]+inp_5[53];
  assign {FA_cout_118,FA_out_118}=inp_3[56]+inp_4[55]+inp_5[54];
  assign {FA_cout_119,FA_out_119}=inp_3[57]+inp_4[56]+inp_5[55];
  assign {FA_cout_120,FA_out_120}=inp_3[58]+inp_4[57]+inp_5[56];
  assign {FA_cout_121,FA_out_121}=inp_3[59]+inp_4[58]+inp_5[57];
  assign {FA_cout_122,FA_out_122}=inp_3[60]+inp_4[59]+inp_5[58];
  assign {FA_cout_123,FA_out_123}=inp_3[61]+inp_4[60]+inp_5[59];
  assign {FA_cout_124,FA_out_124}=inp_3[63]+inp_4[62]+inp_5[61];
  assign {FA_cout_125,FA_out_125}=inp_4[63]+inp_5[62]+inp_6[61];
  assign {FA_cout_126,FA_out_126}=inp_5[60]+inp_6[59]+inp_7[58];
  assign {FA_cout_127,FA_out_127}=inp_5[63]+inp_6[62]+inp_7[61];
  assign {FA_cout_128,FA_out_128}=inp_6[2]+inp_7[1]+inp_8[0];
  assign {FA_cout_129,FA_out_129}=inp_6[3]+inp_7[2]+inp_8[1];
  assign {FA_cout_130,FA_out_130}=inp_6[4]+inp_7[3]+inp_8[2];
  assign {FA_cout_131,FA_out_131}=inp_6[5]+inp_7[4]+inp_8[3];
  assign {FA_cout_132,FA_out_132}=inp_6[6]+inp_7[5]+inp_8[4];
  assign {FA_cout_133,FA_out_133}=inp_6[7]+inp_7[6]+inp_8[5];
  assign {FA_cout_134,FA_out_134}=inp_6[8]+inp_7[7]+inp_8[6];
  assign {FA_cout_135,FA_out_135}=inp_6[9]+inp_7[8]+inp_8[7];
  assign {FA_cout_136,FA_out_136}=inp_6[10]+inp_7[9]+inp_8[8];
  assign {FA_cout_137,FA_out_137}=inp_6[11]+inp_7[10]+inp_8[9];
  assign {FA_cout_138,FA_out_138}=inp_6[12]+inp_7[11]+inp_8[10];
  assign {FA_cout_139,FA_out_139}=inp_6[13]+inp_7[12]+inp_8[11];
  assign {FA_cout_140,FA_out_140}=inp_6[14]+inp_7[13]+inp_8[12];
  assign {FA_cout_141,FA_out_141}=inp_6[15]+inp_7[14]+inp_8[13];
  assign {FA_cout_142,FA_out_142}=inp_6[16]+inp_7[15]+inp_8[14];
  assign {FA_cout_143,FA_out_143}=inp_6[17]+inp_7[16]+inp_8[15];
  assign {FA_cout_144,FA_out_144}=inp_6[18]+inp_7[17]+inp_8[16];
  assign {FA_cout_145,FA_out_145}=inp_6[19]+inp_7[18]+inp_8[17];
  assign {FA_cout_146,FA_out_146}=inp_6[20]+inp_7[19]+inp_8[18];
  assign {FA_cout_147,FA_out_147}=inp_6[21]+inp_7[20]+inp_8[19];
  assign {FA_cout_148,FA_out_148}=inp_6[22]+inp_7[21]+inp_8[20];
  assign {FA_cout_149,FA_out_149}=inp_6[23]+inp_7[22]+inp_8[21];
  assign {FA_cout_150,FA_out_150}=inp_6[24]+inp_7[23]+inp_8[22];
  assign {FA_cout_151,FA_out_151}=inp_6[25]+inp_7[24]+inp_8[23];
  assign {FA_cout_152,FA_out_152}=inp_6[26]+inp_7[25]+inp_8[24];
  assign {FA_cout_153,FA_out_153}=inp_6[27]+inp_7[26]+inp_8[25];
  assign {FA_cout_154,FA_out_154}=inp_6[28]+inp_7[27]+inp_8[26];
  assign {FA_cout_155,FA_out_155}=inp_6[29]+inp_7[28]+inp_8[27];
  assign {FA_cout_156,FA_out_156}=inp_6[30]+inp_7[29]+inp_8[28];
  assign {FA_cout_157,FA_out_157}=inp_6[31]+inp_7[30]+inp_8[29];
  assign {FA_cout_158,FA_out_158}=inp_6[32]+inp_7[31]+inp_8[30];
  assign {FA_cout_159,FA_out_159}=inp_6[33]+inp_7[32]+inp_8[31];
  assign {FA_cout_160,FA_out_160}=inp_6[34]+inp_7[33]+inp_8[32];
  assign {FA_cout_161,FA_out_161}=inp_6[35]+inp_7[34]+inp_8[33];
  assign {FA_cout_162,FA_out_162}=inp_6[36]+inp_7[35]+inp_8[34];
  assign {FA_cout_163,FA_out_163}=inp_6[37]+inp_7[36]+inp_8[35];
  assign {FA_cout_164,FA_out_164}=inp_6[38]+inp_7[37]+inp_8[36];
  assign {FA_cout_165,FA_out_165}=inp_6[39]+inp_7[38]+inp_8[37];
  assign {FA_cout_166,FA_out_166}=inp_6[40]+inp_7[39]+inp_8[38];
  assign {FA_cout_167,FA_out_167}=inp_6[41]+inp_7[40]+inp_8[39];
  assign {FA_cout_168,FA_out_168}=inp_6[42]+inp_7[41]+inp_8[40];
  assign {FA_cout_169,FA_out_169}=inp_6[43]+inp_7[42]+inp_8[41];
  assign {FA_cout_170,FA_out_170}=inp_6[44]+inp_7[43]+inp_8[42];
  assign {FA_cout_171,FA_out_171}=inp_6[45]+inp_7[44]+inp_8[43];
  assign {FA_cout_172,FA_out_172}=inp_6[46]+inp_7[45]+inp_8[44];
  assign {FA_cout_173,FA_out_173}=inp_6[47]+inp_7[46]+inp_8[45];
  assign {FA_cout_174,FA_out_174}=inp_6[48]+inp_7[47]+inp_8[46];
  assign {FA_cout_175,FA_out_175}=inp_6[49]+inp_7[48]+inp_8[47];
  assign {FA_cout_176,FA_out_176}=inp_6[50]+inp_7[49]+inp_8[48];
  assign {FA_cout_177,FA_out_177}=inp_6[51]+inp_7[50]+inp_8[49];
  assign {FA_cout_178,FA_out_178}=inp_6[52]+inp_7[51]+inp_8[50];
  assign {FA_cout_179,FA_out_179}=inp_6[53]+inp_7[52]+inp_8[51];
  assign {FA_cout_180,FA_out_180}=inp_6[54]+inp_7[53]+inp_8[52];
  assign {FA_cout_181,FA_out_181}=inp_6[55]+inp_7[54]+inp_8[53];
  assign {FA_cout_182,FA_out_182}=inp_6[56]+inp_7[55]+inp_8[54];
  assign {FA_cout_183,FA_out_183}=inp_6[57]+inp_7[56]+inp_8[55];
  assign {FA_cout_184,FA_out_184}=inp_6[58]+inp_7[57]+inp_8[56];
  assign {FA_cout_185,FA_out_185}=inp_6[60]+inp_7[59]+inp_8[58];
  assign {FA_cout_186,FA_out_186}=inp_6[63]+inp_7[62]+inp_8[61];
  assign {FA_cout_187,FA_out_187}=inp_7[60]+inp_8[59]+inp_9[58];
  assign {FA_cout_188,FA_out_188}=inp_7[63]+inp_8[62]+inp_9[61];
  assign {FA_cout_189,FA_out_189}=inp_8[57]+inp_9[56]+inp_10[55];
  assign {FA_cout_190,FA_out_190}=inp_8[60]+inp_9[59]+inp_10[58];
  assign {FA_cout_191,FA_out_191}=inp_8[63]+inp_9[62]+inp_10[61];
  assign {FA_cout_192,FA_out_192}=inp_9[2]+inp_10[1]+inp_11[0];
  assign {FA_cout_193,FA_out_193}=inp_9[3]+inp_10[2]+inp_11[1];
  assign {FA_cout_194,FA_out_194}=inp_9[4]+inp_10[3]+inp_11[2];
  assign {FA_cout_195,FA_out_195}=inp_9[5]+inp_10[4]+inp_11[3];
  assign {FA_cout_196,FA_out_196}=inp_9[6]+inp_10[5]+inp_11[4];
  assign {FA_cout_197,FA_out_197}=inp_9[7]+inp_10[6]+inp_11[5];
  assign {FA_cout_198,FA_out_198}=inp_9[8]+inp_10[7]+inp_11[6];
  assign {FA_cout_199,FA_out_199}=inp_9[9]+inp_10[8]+inp_11[7];
  assign {FA_cout_200,FA_out_200}=inp_9[10]+inp_10[9]+inp_11[8];
  assign {FA_cout_201,FA_out_201}=inp_9[11]+inp_10[10]+inp_11[9];
  assign {FA_cout_202,FA_out_202}=inp_9[12]+inp_10[11]+inp_11[10];
  assign {FA_cout_203,FA_out_203}=inp_9[13]+inp_10[12]+inp_11[11];
  assign {FA_cout_204,FA_out_204}=inp_9[14]+inp_10[13]+inp_11[12];
  assign {FA_cout_205,FA_out_205}=inp_9[15]+inp_10[14]+inp_11[13];
  assign {FA_cout_206,FA_out_206}=inp_9[16]+inp_10[15]+inp_11[14];
  assign {FA_cout_207,FA_out_207}=inp_9[17]+inp_10[16]+inp_11[15];
  assign {FA_cout_208,FA_out_208}=inp_9[18]+inp_10[17]+inp_11[16];
  assign {FA_cout_209,FA_out_209}=inp_9[19]+inp_10[18]+inp_11[17];
  assign {FA_cout_210,FA_out_210}=inp_9[20]+inp_10[19]+inp_11[18];
  assign {FA_cout_211,FA_out_211}=inp_9[21]+inp_10[20]+inp_11[19];
  assign {FA_cout_212,FA_out_212}=inp_9[22]+inp_10[21]+inp_11[20];
  assign {FA_cout_213,FA_out_213}=inp_9[23]+inp_10[22]+inp_11[21];
  assign {FA_cout_214,FA_out_214}=inp_9[24]+inp_10[23]+inp_11[22];
  assign {FA_cout_215,FA_out_215}=inp_9[25]+inp_10[24]+inp_11[23];
  assign {FA_cout_216,FA_out_216}=inp_9[26]+inp_10[25]+inp_11[24];
  assign {FA_cout_217,FA_out_217}=inp_9[27]+inp_10[26]+inp_11[25];
  assign {FA_cout_218,FA_out_218}=inp_9[28]+inp_10[27]+inp_11[26];
  assign {FA_cout_219,FA_out_219}=inp_9[29]+inp_10[28]+inp_11[27];
  assign {FA_cout_220,FA_out_220}=inp_9[30]+inp_10[29]+inp_11[28];
  assign {FA_cout_221,FA_out_221}=inp_9[31]+inp_10[30]+inp_11[29];
  assign {FA_cout_222,FA_out_222}=inp_9[32]+inp_10[31]+inp_11[30];
  assign {FA_cout_223,FA_out_223}=inp_9[33]+inp_10[32]+inp_11[31];
  assign {FA_cout_224,FA_out_224}=inp_9[34]+inp_10[33]+inp_11[32];
  assign {FA_cout_225,FA_out_225}=inp_9[35]+inp_10[34]+inp_11[33];
  assign {FA_cout_226,FA_out_226}=inp_9[36]+inp_10[35]+inp_11[34];
  assign {FA_cout_227,FA_out_227}=inp_9[37]+inp_10[36]+inp_11[35];
  assign {FA_cout_228,FA_out_228}=inp_9[38]+inp_10[37]+inp_11[36];
  assign {FA_cout_229,FA_out_229}=inp_9[39]+inp_10[38]+inp_11[37];
  assign {FA_cout_230,FA_out_230}=inp_9[40]+inp_10[39]+inp_11[38];
  assign {FA_cout_231,FA_out_231}=inp_9[41]+inp_10[40]+inp_11[39];
  assign {FA_cout_232,FA_out_232}=inp_9[42]+inp_10[41]+inp_11[40];
  assign {FA_cout_233,FA_out_233}=inp_9[43]+inp_10[42]+inp_11[41];
  assign {FA_cout_234,FA_out_234}=inp_9[44]+inp_10[43]+inp_11[42];
  assign {FA_cout_235,FA_out_235}=inp_9[45]+inp_10[44]+inp_11[43];
  assign {FA_cout_236,FA_out_236}=inp_9[46]+inp_10[45]+inp_11[44];
  assign {FA_cout_237,FA_out_237}=inp_9[47]+inp_10[46]+inp_11[45];
  assign {FA_cout_238,FA_out_238}=inp_9[48]+inp_10[47]+inp_11[46];
  assign {FA_cout_239,FA_out_239}=inp_9[49]+inp_10[48]+inp_11[47];
  assign {FA_cout_240,FA_out_240}=inp_9[50]+inp_10[49]+inp_11[48];
  assign {FA_cout_241,FA_out_241}=inp_9[51]+inp_10[50]+inp_11[49];
  assign {FA_cout_242,FA_out_242}=inp_9[52]+inp_10[51]+inp_11[50];
  assign {FA_cout_243,FA_out_243}=inp_9[53]+inp_10[52]+inp_11[51];
  assign {FA_cout_244,FA_out_244}=inp_9[54]+inp_10[53]+inp_11[52];
  assign {FA_cout_245,FA_out_245}=inp_9[55]+inp_10[54]+inp_11[53];
  assign {FA_cout_246,FA_out_246}=inp_9[57]+inp_10[56]+inp_11[55];
  assign {FA_cout_247,FA_out_247}=inp_9[60]+inp_10[59]+inp_11[58];
  assign {FA_cout_248,FA_out_248}=inp_9[63]+inp_10[62]+inp_11[61];
  assign {FA_cout_249,FA_out_249}=inp_10[57]+inp_11[56]+inp_12[55];
  assign {FA_cout_250,FA_out_250}=inp_10[60]+inp_11[59]+inp_12[58];
  assign {FA_cout_251,FA_out_251}=inp_10[63]+inp_11[62]+inp_12[61];
  assign {FA_cout_252,FA_out_252}=inp_11[54]+inp_12[53]+inp_13[52];
  assign {FA_cout_253,FA_out_253}=inp_11[57]+inp_12[56]+inp_13[55];
  assign {FA_cout_254,FA_out_254}=inp_11[60]+inp_12[59]+inp_13[58];
  assign {FA_cout_255,FA_out_255}=inp_11[63]+inp_12[62]+inp_13[61];
  assign {FA_cout_256,FA_out_256}=inp_12[2]+inp_13[1]+inp_14[0];
  assign {FA_cout_257,FA_out_257}=inp_12[3]+inp_13[2]+inp_14[1];
  assign {FA_cout_258,FA_out_258}=inp_12[4]+inp_13[3]+inp_14[2];
  assign {FA_cout_259,FA_out_259}=inp_12[5]+inp_13[4]+inp_14[3];
  assign {FA_cout_260,FA_out_260}=inp_12[6]+inp_13[5]+inp_14[4];
  assign {FA_cout_261,FA_out_261}=inp_12[7]+inp_13[6]+inp_14[5];
  assign {FA_cout_262,FA_out_262}=inp_12[8]+inp_13[7]+inp_14[6];
  assign {FA_cout_263,FA_out_263}=inp_12[9]+inp_13[8]+inp_14[7];
  assign {FA_cout_264,FA_out_264}=inp_12[10]+inp_13[9]+inp_14[8];
  assign {FA_cout_265,FA_out_265}=inp_12[11]+inp_13[10]+inp_14[9];
  assign {FA_cout_266,FA_out_266}=inp_12[12]+inp_13[11]+inp_14[10];
  assign {FA_cout_267,FA_out_267}=inp_12[13]+inp_13[12]+inp_14[11];
  assign {FA_cout_268,FA_out_268}=inp_12[14]+inp_13[13]+inp_14[12];
  assign {FA_cout_269,FA_out_269}=inp_12[15]+inp_13[14]+inp_14[13];
  assign {FA_cout_270,FA_out_270}=inp_12[16]+inp_13[15]+inp_14[14];
  assign {FA_cout_271,FA_out_271}=inp_12[17]+inp_13[16]+inp_14[15];
  assign {FA_cout_272,FA_out_272}=inp_12[18]+inp_13[17]+inp_14[16];
  assign {FA_cout_273,FA_out_273}=inp_12[19]+inp_13[18]+inp_14[17];
  assign {FA_cout_274,FA_out_274}=inp_12[20]+inp_13[19]+inp_14[18];
  assign {FA_cout_275,FA_out_275}=inp_12[21]+inp_13[20]+inp_14[19];
  assign {FA_cout_276,FA_out_276}=inp_12[22]+inp_13[21]+inp_14[20];
  assign {FA_cout_277,FA_out_277}=inp_12[23]+inp_13[22]+inp_14[21];
  assign {FA_cout_278,FA_out_278}=inp_12[24]+inp_13[23]+inp_14[22];
  assign {FA_cout_279,FA_out_279}=inp_12[25]+inp_13[24]+inp_14[23];
  assign {FA_cout_280,FA_out_280}=inp_12[26]+inp_13[25]+inp_14[24];
  assign {FA_cout_281,FA_out_281}=inp_12[27]+inp_13[26]+inp_14[25];
  assign {FA_cout_282,FA_out_282}=inp_12[28]+inp_13[27]+inp_14[26];
  assign {FA_cout_283,FA_out_283}=inp_12[29]+inp_13[28]+inp_14[27];
  assign {FA_cout_284,FA_out_284}=inp_12[30]+inp_13[29]+inp_14[28];
  assign {FA_cout_285,FA_out_285}=inp_12[31]+inp_13[30]+inp_14[29];
  assign {FA_cout_286,FA_out_286}=inp_12[32]+inp_13[31]+inp_14[30];
  assign {FA_cout_287,FA_out_287}=inp_12[33]+inp_13[32]+inp_14[31];
  assign {FA_cout_288,FA_out_288}=inp_12[34]+inp_13[33]+inp_14[32];
  assign {FA_cout_289,FA_out_289}=inp_12[35]+inp_13[34]+inp_14[33];
  assign {FA_cout_290,FA_out_290}=inp_12[36]+inp_13[35]+inp_14[34];
  assign {FA_cout_291,FA_out_291}=inp_12[37]+inp_13[36]+inp_14[35];
  assign {FA_cout_292,FA_out_292}=inp_12[38]+inp_13[37]+inp_14[36];
  assign {FA_cout_293,FA_out_293}=inp_12[39]+inp_13[38]+inp_14[37];
  assign {FA_cout_294,FA_out_294}=inp_12[40]+inp_13[39]+inp_14[38];
  assign {FA_cout_295,FA_out_295}=inp_12[41]+inp_13[40]+inp_14[39];
  assign {FA_cout_296,FA_out_296}=inp_12[42]+inp_13[41]+inp_14[40];
  assign {FA_cout_297,FA_out_297}=inp_12[43]+inp_13[42]+inp_14[41];
  assign {FA_cout_298,FA_out_298}=inp_12[44]+inp_13[43]+inp_14[42];
  assign {FA_cout_299,FA_out_299}=inp_12[45]+inp_13[44]+inp_14[43];
  assign {FA_cout_300,FA_out_300}=inp_12[46]+inp_13[45]+inp_14[44];
  assign {FA_cout_301,FA_out_301}=inp_12[47]+inp_13[46]+inp_14[45];
  assign {FA_cout_302,FA_out_302}=inp_12[48]+inp_13[47]+inp_14[46];
  assign {FA_cout_303,FA_out_303}=inp_12[49]+inp_13[48]+inp_14[47];
  assign {FA_cout_304,FA_out_304}=inp_12[50]+inp_13[49]+inp_14[48];
  assign {FA_cout_305,FA_out_305}=inp_12[51]+inp_13[50]+inp_14[49];
  assign {FA_cout_306,FA_out_306}=inp_12[52]+inp_13[51]+inp_14[50];
  assign {FA_cout_307,FA_out_307}=inp_12[54]+inp_13[53]+inp_14[52];
  assign {FA_cout_308,FA_out_308}=inp_12[57]+inp_13[56]+inp_14[55];
  assign {FA_cout_309,FA_out_309}=inp_12[60]+inp_13[59]+inp_14[58];
  assign {FA_cout_310,FA_out_310}=inp_12[63]+inp_13[62]+inp_14[61];
  assign {FA_cout_311,FA_out_311}=inp_13[54]+inp_14[53]+inp_15[52];
  assign {FA_cout_312,FA_out_312}=inp_13[57]+inp_14[56]+inp_15[55];
  assign {FA_cout_313,FA_out_313}=inp_13[60]+inp_14[59]+inp_15[58];
  assign {FA_cout_314,FA_out_314}=inp_13[63]+inp_14[62]+inp_15[61];
  assign {FA_cout_315,FA_out_315}=inp_14[51]+inp_15[50]+inp_16[49];
  assign {FA_cout_316,FA_out_316}=inp_14[54]+inp_15[53]+inp_16[52];
  assign {FA_cout_317,FA_out_317}=inp_14[57]+inp_15[56]+inp_16[55];
  assign {FA_cout_318,FA_out_318}=inp_14[60]+inp_15[59]+inp_16[58];
  assign {FA_cout_319,FA_out_319}=inp_14[63]+inp_15[62]+inp_16[61];
  assign {FA_cout_320,FA_out_320}=inp_15[2]+inp_16[1]+inp_17[0];
  assign {FA_cout_321,FA_out_321}=inp_15[3]+inp_16[2]+inp_17[1];
  assign {FA_cout_322,FA_out_322}=inp_15[4]+inp_16[3]+inp_17[2];
  assign {FA_cout_323,FA_out_323}=inp_15[5]+inp_16[4]+inp_17[3];
  assign {FA_cout_324,FA_out_324}=inp_15[6]+inp_16[5]+inp_17[4];
  assign {FA_cout_325,FA_out_325}=inp_15[7]+inp_16[6]+inp_17[5];
  assign {FA_cout_326,FA_out_326}=inp_15[8]+inp_16[7]+inp_17[6];
  assign {FA_cout_327,FA_out_327}=inp_15[9]+inp_16[8]+inp_17[7];
  assign {FA_cout_328,FA_out_328}=inp_15[10]+inp_16[9]+inp_17[8];
  assign {FA_cout_329,FA_out_329}=inp_15[11]+inp_16[10]+inp_17[9];
  assign {FA_cout_330,FA_out_330}=inp_15[12]+inp_16[11]+inp_17[10];
  assign {FA_cout_331,FA_out_331}=inp_15[13]+inp_16[12]+inp_17[11];
  assign {FA_cout_332,FA_out_332}=inp_15[14]+inp_16[13]+inp_17[12];
  assign {FA_cout_333,FA_out_333}=inp_15[15]+inp_16[14]+inp_17[13];
  assign {FA_cout_334,FA_out_334}=inp_15[16]+inp_16[15]+inp_17[14];
  assign {FA_cout_335,FA_out_335}=inp_15[17]+inp_16[16]+inp_17[15];
  assign {FA_cout_336,FA_out_336}=inp_15[18]+inp_16[17]+inp_17[16];
  assign {FA_cout_337,FA_out_337}=inp_15[19]+inp_16[18]+inp_17[17];
  assign {FA_cout_338,FA_out_338}=inp_15[20]+inp_16[19]+inp_17[18];
  assign {FA_cout_339,FA_out_339}=inp_15[21]+inp_16[20]+inp_17[19];
  assign {FA_cout_340,FA_out_340}=inp_15[22]+inp_16[21]+inp_17[20];
  assign {FA_cout_341,FA_out_341}=inp_15[23]+inp_16[22]+inp_17[21];
  assign {FA_cout_342,FA_out_342}=inp_15[24]+inp_16[23]+inp_17[22];
  assign {FA_cout_343,FA_out_343}=inp_15[25]+inp_16[24]+inp_17[23];
  assign {FA_cout_344,FA_out_344}=inp_15[26]+inp_16[25]+inp_17[24];
  assign {FA_cout_345,FA_out_345}=inp_15[27]+inp_16[26]+inp_17[25];
  assign {FA_cout_346,FA_out_346}=inp_15[28]+inp_16[27]+inp_17[26];
  assign {FA_cout_347,FA_out_347}=inp_15[29]+inp_16[28]+inp_17[27];
  assign {FA_cout_348,FA_out_348}=inp_15[30]+inp_16[29]+inp_17[28];
  assign {FA_cout_349,FA_out_349}=inp_15[31]+inp_16[30]+inp_17[29];
  assign {FA_cout_350,FA_out_350}=inp_15[32]+inp_16[31]+inp_17[30];
  assign {FA_cout_351,FA_out_351}=inp_15[33]+inp_16[32]+inp_17[31];
  assign {FA_cout_352,FA_out_352}=inp_15[34]+inp_16[33]+inp_17[32];
  assign {FA_cout_353,FA_out_353}=inp_15[35]+inp_16[34]+inp_17[33];
  assign {FA_cout_354,FA_out_354}=inp_15[36]+inp_16[35]+inp_17[34];
  assign {FA_cout_355,FA_out_355}=inp_15[37]+inp_16[36]+inp_17[35];
  assign {FA_cout_356,FA_out_356}=inp_15[38]+inp_16[37]+inp_17[36];
  assign {FA_cout_357,FA_out_357}=inp_15[39]+inp_16[38]+inp_17[37];
  assign {FA_cout_358,FA_out_358}=inp_15[40]+inp_16[39]+inp_17[38];
  assign {FA_cout_359,FA_out_359}=inp_15[41]+inp_16[40]+inp_17[39];
  assign {FA_cout_360,FA_out_360}=inp_15[42]+inp_16[41]+inp_17[40];
  assign {FA_cout_361,FA_out_361}=inp_15[43]+inp_16[42]+inp_17[41];
  assign {FA_cout_362,FA_out_362}=inp_15[44]+inp_16[43]+inp_17[42];
  assign {FA_cout_363,FA_out_363}=inp_15[45]+inp_16[44]+inp_17[43];
  assign {FA_cout_364,FA_out_364}=inp_15[46]+inp_16[45]+inp_17[44];
  assign {FA_cout_365,FA_out_365}=inp_15[47]+inp_16[46]+inp_17[45];
  assign {FA_cout_366,FA_out_366}=inp_15[48]+inp_16[47]+inp_17[46];
  assign {FA_cout_367,FA_out_367}=inp_15[49]+inp_16[48]+inp_17[47];
  assign {FA_cout_368,FA_out_368}=inp_15[51]+inp_16[50]+inp_17[49];
  assign {FA_cout_369,FA_out_369}=inp_15[54]+inp_16[53]+inp_17[52];
  assign {FA_cout_370,FA_out_370}=inp_15[57]+inp_16[56]+inp_17[55];
  assign {FA_cout_371,FA_out_371}=inp_15[60]+inp_16[59]+inp_17[58];
  assign {FA_cout_372,FA_out_372}=inp_15[63]+inp_16[62]+inp_17[61];
  assign {FA_cout_373,FA_out_373}=inp_16[51]+inp_17[50]+inp_18[49];
  assign {FA_cout_374,FA_out_374}=inp_16[54]+inp_17[53]+inp_18[52];
  assign {FA_cout_375,FA_out_375}=inp_16[57]+inp_17[56]+inp_18[55];
  assign {FA_cout_376,FA_out_376}=inp_16[60]+inp_17[59]+inp_18[58];
  assign {FA_cout_377,FA_out_377}=inp_16[63]+inp_17[62]+inp_18[61];
  assign {FA_cout_378,FA_out_378}=inp_17[48]+inp_18[47]+inp_19[46];
  assign {FA_cout_379,FA_out_379}=inp_17[51]+inp_18[50]+inp_19[49];
  assign {FA_cout_380,FA_out_380}=inp_17[54]+inp_18[53]+inp_19[52];
  assign {FA_cout_381,FA_out_381}=inp_17[57]+inp_18[56]+inp_19[55];
  assign {FA_cout_382,FA_out_382}=inp_17[60]+inp_18[59]+inp_19[58];
  assign {FA_cout_383,FA_out_383}=inp_17[63]+inp_18[62]+inp_19[61];
  assign {FA_cout_384,FA_out_384}=inp_18[2]+inp_19[1]+inp_20[0];
  assign {FA_cout_385,FA_out_385}=inp_18[3]+inp_19[2]+inp_20[1];
  assign {FA_cout_386,FA_out_386}=inp_18[4]+inp_19[3]+inp_20[2];
  assign {FA_cout_387,FA_out_387}=inp_18[5]+inp_19[4]+inp_20[3];
  assign {FA_cout_388,FA_out_388}=inp_18[6]+inp_19[5]+inp_20[4];
  assign {FA_cout_389,FA_out_389}=inp_18[7]+inp_19[6]+inp_20[5];
  assign {FA_cout_390,FA_out_390}=inp_18[8]+inp_19[7]+inp_20[6];
  assign {FA_cout_391,FA_out_391}=inp_18[9]+inp_19[8]+inp_20[7];
  assign {FA_cout_392,FA_out_392}=inp_18[10]+inp_19[9]+inp_20[8];
  assign {FA_cout_393,FA_out_393}=inp_18[11]+inp_19[10]+inp_20[9];
  assign {FA_cout_394,FA_out_394}=inp_18[12]+inp_19[11]+inp_20[10];
  assign {FA_cout_395,FA_out_395}=inp_18[13]+inp_19[12]+inp_20[11];
  assign {FA_cout_396,FA_out_396}=inp_18[14]+inp_19[13]+inp_20[12];
  assign {FA_cout_397,FA_out_397}=inp_18[15]+inp_19[14]+inp_20[13];
  assign {FA_cout_398,FA_out_398}=inp_18[16]+inp_19[15]+inp_20[14];
  assign {FA_cout_399,FA_out_399}=inp_18[17]+inp_19[16]+inp_20[15];
  assign {FA_cout_400,FA_out_400}=inp_18[18]+inp_19[17]+inp_20[16];
  assign {FA_cout_401,FA_out_401}=inp_18[19]+inp_19[18]+inp_20[17];
  assign {FA_cout_402,FA_out_402}=inp_18[20]+inp_19[19]+inp_20[18];
  assign {FA_cout_403,FA_out_403}=inp_18[21]+inp_19[20]+inp_20[19];
  assign {FA_cout_404,FA_out_404}=inp_18[22]+inp_19[21]+inp_20[20];
  assign {FA_cout_405,FA_out_405}=inp_18[23]+inp_19[22]+inp_20[21];
  assign {FA_cout_406,FA_out_406}=inp_18[24]+inp_19[23]+inp_20[22];
  assign {FA_cout_407,FA_out_407}=inp_18[25]+inp_19[24]+inp_20[23];
  assign {FA_cout_408,FA_out_408}=inp_18[26]+inp_19[25]+inp_20[24];
  assign {FA_cout_409,FA_out_409}=inp_18[27]+inp_19[26]+inp_20[25];
  assign {FA_cout_410,FA_out_410}=inp_18[28]+inp_19[27]+inp_20[26];
  assign {FA_cout_411,FA_out_411}=inp_18[29]+inp_19[28]+inp_20[27];
  assign {FA_cout_412,FA_out_412}=inp_18[30]+inp_19[29]+inp_20[28];
  assign {FA_cout_413,FA_out_413}=inp_18[31]+inp_19[30]+inp_20[29];
  assign {FA_cout_414,FA_out_414}=inp_18[32]+inp_19[31]+inp_20[30];
  assign {FA_cout_415,FA_out_415}=inp_18[33]+inp_19[32]+inp_20[31];
  assign {FA_cout_416,FA_out_416}=inp_18[34]+inp_19[33]+inp_20[32];
  assign {FA_cout_417,FA_out_417}=inp_18[35]+inp_19[34]+inp_20[33];
  assign {FA_cout_418,FA_out_418}=inp_18[36]+inp_19[35]+inp_20[34];
  assign {FA_cout_419,FA_out_419}=inp_18[37]+inp_19[36]+inp_20[35];
  assign {FA_cout_420,FA_out_420}=inp_18[38]+inp_19[37]+inp_20[36];
  assign {FA_cout_421,FA_out_421}=inp_18[39]+inp_19[38]+inp_20[37];
  assign {FA_cout_422,FA_out_422}=inp_18[40]+inp_19[39]+inp_20[38];
  assign {FA_cout_423,FA_out_423}=inp_18[41]+inp_19[40]+inp_20[39];
  assign {FA_cout_424,FA_out_424}=inp_18[42]+inp_19[41]+inp_20[40];
  assign {FA_cout_425,FA_out_425}=inp_18[43]+inp_19[42]+inp_20[41];
  assign {FA_cout_426,FA_out_426}=inp_18[44]+inp_19[43]+inp_20[42];
  assign {FA_cout_427,FA_out_427}=inp_18[45]+inp_19[44]+inp_20[43];
  assign {FA_cout_428,FA_out_428}=inp_18[46]+inp_19[45]+inp_20[44];
  assign {FA_cout_429,FA_out_429}=inp_18[48]+inp_19[47]+inp_20[46];
  assign {FA_cout_430,FA_out_430}=inp_18[51]+inp_19[50]+inp_20[49];
  assign {FA_cout_431,FA_out_431}=inp_18[54]+inp_19[53]+inp_20[52];
  assign {FA_cout_432,FA_out_432}=inp_18[57]+inp_19[56]+inp_20[55];
  assign {FA_cout_433,FA_out_433}=inp_18[60]+inp_19[59]+inp_20[58];
  assign {FA_cout_434,FA_out_434}=inp_18[63]+inp_19[62]+inp_20[61];
  assign {FA_cout_435,FA_out_435}=inp_19[48]+inp_20[47]+inp_21[46];
  assign {FA_cout_436,FA_out_436}=inp_19[51]+inp_20[50]+inp_21[49];
  assign {FA_cout_437,FA_out_437}=inp_19[54]+inp_20[53]+inp_21[52];
  assign {FA_cout_438,FA_out_438}=inp_19[57]+inp_20[56]+inp_21[55];
  assign {FA_cout_439,FA_out_439}=inp_19[60]+inp_20[59]+inp_21[58];
  assign {FA_cout_440,FA_out_440}=inp_19[63]+inp_20[62]+inp_21[61];
  assign {FA_cout_441,FA_out_441}=inp_20[45]+inp_21[44]+inp_22[43];
  assign {FA_cout_442,FA_out_442}=inp_20[48]+inp_21[47]+inp_22[46];
  assign {FA_cout_443,FA_out_443}=inp_20[51]+inp_21[50]+inp_22[49];
  assign {FA_cout_444,FA_out_444}=inp_20[54]+inp_21[53]+inp_22[52];
  assign {FA_cout_445,FA_out_445}=inp_20[57]+inp_21[56]+inp_22[55];
  assign {FA_cout_446,FA_out_446}=inp_20[60]+inp_21[59]+inp_22[58];
  assign {FA_cout_447,FA_out_447}=inp_20[63]+inp_21[62]+inp_22[61];
  assign {FA_cout_448,FA_out_448}=inp_21[2]+inp_22[1]+inp_23[0];
  assign {FA_cout_449,FA_out_449}=inp_21[3]+inp_22[2]+inp_23[1];
  assign {FA_cout_450,FA_out_450}=inp_21[4]+inp_22[3]+inp_23[2];
  assign {FA_cout_451,FA_out_451}=inp_21[5]+inp_22[4]+inp_23[3];
  assign {FA_cout_452,FA_out_452}=inp_21[6]+inp_22[5]+inp_23[4];
  assign {FA_cout_453,FA_out_453}=inp_21[7]+inp_22[6]+inp_23[5];
  assign {FA_cout_454,FA_out_454}=inp_21[8]+inp_22[7]+inp_23[6];
  assign {FA_cout_455,FA_out_455}=inp_21[9]+inp_22[8]+inp_23[7];
  assign {FA_cout_456,FA_out_456}=inp_21[10]+inp_22[9]+inp_23[8];
  assign {FA_cout_457,FA_out_457}=inp_21[11]+inp_22[10]+inp_23[9];
  assign {FA_cout_458,FA_out_458}=inp_21[12]+inp_22[11]+inp_23[10];
  assign {FA_cout_459,FA_out_459}=inp_21[13]+inp_22[12]+inp_23[11];
  assign {FA_cout_460,FA_out_460}=inp_21[14]+inp_22[13]+inp_23[12];
  assign {FA_cout_461,FA_out_461}=inp_21[15]+inp_22[14]+inp_23[13];
  assign {FA_cout_462,FA_out_462}=inp_21[16]+inp_22[15]+inp_23[14];
  assign {FA_cout_463,FA_out_463}=inp_21[17]+inp_22[16]+inp_23[15];
  assign {FA_cout_464,FA_out_464}=inp_21[18]+inp_22[17]+inp_23[16];
  assign {FA_cout_465,FA_out_465}=inp_21[19]+inp_22[18]+inp_23[17];
  assign {FA_cout_466,FA_out_466}=inp_21[20]+inp_22[19]+inp_23[18];
  assign {FA_cout_467,FA_out_467}=inp_21[21]+inp_22[20]+inp_23[19];
  assign {FA_cout_468,FA_out_468}=inp_21[22]+inp_22[21]+inp_23[20];
  assign {FA_cout_469,FA_out_469}=inp_21[23]+inp_22[22]+inp_23[21];
  assign {FA_cout_470,FA_out_470}=inp_21[24]+inp_22[23]+inp_23[22];
  assign {FA_cout_471,FA_out_471}=inp_21[25]+inp_22[24]+inp_23[23];
  assign {FA_cout_472,FA_out_472}=inp_21[26]+inp_22[25]+inp_23[24];
  assign {FA_cout_473,FA_out_473}=inp_21[27]+inp_22[26]+inp_23[25];
  assign {FA_cout_474,FA_out_474}=inp_21[28]+inp_22[27]+inp_23[26];
  assign {FA_cout_475,FA_out_475}=inp_21[29]+inp_22[28]+inp_23[27];
  assign {FA_cout_476,FA_out_476}=inp_21[30]+inp_22[29]+inp_23[28];
  assign {FA_cout_477,FA_out_477}=inp_21[31]+inp_22[30]+inp_23[29];
  assign {FA_cout_478,FA_out_478}=inp_21[32]+inp_22[31]+inp_23[30];
  assign {FA_cout_479,FA_out_479}=inp_21[33]+inp_22[32]+inp_23[31];
  assign {FA_cout_480,FA_out_480}=inp_21[34]+inp_22[33]+inp_23[32];
  assign {FA_cout_481,FA_out_481}=inp_21[35]+inp_22[34]+inp_23[33];
  assign {FA_cout_482,FA_out_482}=inp_21[36]+inp_22[35]+inp_23[34];
  assign {FA_cout_483,FA_out_483}=inp_21[37]+inp_22[36]+inp_23[35];
  assign {FA_cout_484,FA_out_484}=inp_21[38]+inp_22[37]+inp_23[36];
  assign {FA_cout_485,FA_out_485}=inp_21[39]+inp_22[38]+inp_23[37];
  assign {FA_cout_486,FA_out_486}=inp_21[40]+inp_22[39]+inp_23[38];
  assign {FA_cout_487,FA_out_487}=inp_21[41]+inp_22[40]+inp_23[39];
  assign {FA_cout_488,FA_out_488}=inp_21[42]+inp_22[41]+inp_23[40];
  assign {FA_cout_489,FA_out_489}=inp_21[43]+inp_22[42]+inp_23[41];
  assign {FA_cout_490,FA_out_490}=inp_21[45]+inp_22[44]+inp_23[43];
  assign {FA_cout_491,FA_out_491}=inp_21[48]+inp_22[47]+inp_23[46];
  assign {FA_cout_492,FA_out_492}=inp_21[51]+inp_22[50]+inp_23[49];
  assign {FA_cout_493,FA_out_493}=inp_21[54]+inp_22[53]+inp_23[52];
  assign {FA_cout_494,FA_out_494}=inp_21[57]+inp_22[56]+inp_23[55];
  assign {FA_cout_495,FA_out_495}=inp_21[60]+inp_22[59]+inp_23[58];
  assign {FA_cout_496,FA_out_496}=inp_21[63]+inp_22[62]+inp_23[61];
  assign {FA_cout_497,FA_out_497}=inp_22[45]+inp_23[44]+inp_24[43];
  assign {FA_cout_498,FA_out_498}=inp_22[48]+inp_23[47]+inp_24[46];
  assign {FA_cout_499,FA_out_499}=inp_22[51]+inp_23[50]+inp_24[49];
  assign {FA_cout_500,FA_out_500}=inp_22[54]+inp_23[53]+inp_24[52];
  assign {FA_cout_501,FA_out_501}=inp_22[57]+inp_23[56]+inp_24[55];
  assign {FA_cout_502,FA_out_502}=inp_22[60]+inp_23[59]+inp_24[58];
  assign {FA_cout_503,FA_out_503}=inp_22[63]+inp_23[62]+inp_24[61];
  assign {FA_cout_504,FA_out_504}=inp_23[42]+inp_24[41]+inp_25[40];
  assign {FA_cout_505,FA_out_505}=inp_23[45]+inp_24[44]+inp_25[43];
  assign {FA_cout_506,FA_out_506}=inp_23[48]+inp_24[47]+inp_25[46];
  assign {FA_cout_507,FA_out_507}=inp_23[51]+inp_24[50]+inp_25[49];
  assign {FA_cout_508,FA_out_508}=inp_23[54]+inp_24[53]+inp_25[52];
  assign {FA_cout_509,FA_out_509}=inp_23[57]+inp_24[56]+inp_25[55];
  assign {FA_cout_510,FA_out_510}=inp_23[60]+inp_24[59]+inp_25[58];
  assign {FA_cout_511,FA_out_511}=inp_23[63]+inp_24[62]+inp_25[61];
  assign {FA_cout_512,FA_out_512}=inp_24[2]+inp_25[1]+inp_26[0];
  assign {FA_cout_513,FA_out_513}=inp_24[3]+inp_25[2]+inp_26[1];
  assign {FA_cout_514,FA_out_514}=inp_24[4]+inp_25[3]+inp_26[2];
  assign {FA_cout_515,FA_out_515}=inp_24[5]+inp_25[4]+inp_26[3];
  assign {FA_cout_516,FA_out_516}=inp_24[6]+inp_25[5]+inp_26[4];
  assign {FA_cout_517,FA_out_517}=inp_24[7]+inp_25[6]+inp_26[5];
  assign {FA_cout_518,FA_out_518}=inp_24[8]+inp_25[7]+inp_26[6];
  assign {FA_cout_519,FA_out_519}=inp_24[9]+inp_25[8]+inp_26[7];
  assign {FA_cout_520,FA_out_520}=inp_24[10]+inp_25[9]+inp_26[8];
  assign {FA_cout_521,FA_out_521}=inp_24[11]+inp_25[10]+inp_26[9];
  assign {FA_cout_522,FA_out_522}=inp_24[12]+inp_25[11]+inp_26[10];
  assign {FA_cout_523,FA_out_523}=inp_24[13]+inp_25[12]+inp_26[11];
  assign {FA_cout_524,FA_out_524}=inp_24[14]+inp_25[13]+inp_26[12];
  assign {FA_cout_525,FA_out_525}=inp_24[15]+inp_25[14]+inp_26[13];
  assign {FA_cout_526,FA_out_526}=inp_24[16]+inp_25[15]+inp_26[14];
  assign {FA_cout_527,FA_out_527}=inp_24[17]+inp_25[16]+inp_26[15];
  assign {FA_cout_528,FA_out_528}=inp_24[18]+inp_25[17]+inp_26[16];
  assign {FA_cout_529,FA_out_529}=inp_24[19]+inp_25[18]+inp_26[17];
  assign {FA_cout_530,FA_out_530}=inp_24[20]+inp_25[19]+inp_26[18];
  assign {FA_cout_531,FA_out_531}=inp_24[21]+inp_25[20]+inp_26[19];
  assign {FA_cout_532,FA_out_532}=inp_24[22]+inp_25[21]+inp_26[20];
  assign {FA_cout_533,FA_out_533}=inp_24[23]+inp_25[22]+inp_26[21];
  assign {FA_cout_534,FA_out_534}=inp_24[24]+inp_25[23]+inp_26[22];
  assign {FA_cout_535,FA_out_535}=inp_24[25]+inp_25[24]+inp_26[23];
  assign {FA_cout_536,FA_out_536}=inp_24[26]+inp_25[25]+inp_26[24];
  assign {FA_cout_537,FA_out_537}=inp_24[27]+inp_25[26]+inp_26[25];
  assign {FA_cout_538,FA_out_538}=inp_24[28]+inp_25[27]+inp_26[26];
  assign {FA_cout_539,FA_out_539}=inp_24[29]+inp_25[28]+inp_26[27];
  assign {FA_cout_540,FA_out_540}=inp_24[30]+inp_25[29]+inp_26[28];
  assign {FA_cout_541,FA_out_541}=inp_24[31]+inp_25[30]+inp_26[29];
  assign {FA_cout_542,FA_out_542}=inp_24[32]+inp_25[31]+inp_26[30];
  assign {FA_cout_543,FA_out_543}=inp_24[33]+inp_25[32]+inp_26[31];
  assign {FA_cout_544,FA_out_544}=inp_24[34]+inp_25[33]+inp_26[32];
  assign {FA_cout_545,FA_out_545}=inp_24[35]+inp_25[34]+inp_26[33];
  assign {FA_cout_546,FA_out_546}=inp_24[36]+inp_25[35]+inp_26[34];
  assign {FA_cout_547,FA_out_547}=inp_24[37]+inp_25[36]+inp_26[35];
  assign {FA_cout_548,FA_out_548}=inp_24[38]+inp_25[37]+inp_26[36];
  assign {FA_cout_549,FA_out_549}=inp_24[39]+inp_25[38]+inp_26[37];
  assign {FA_cout_550,FA_out_550}=inp_24[40]+inp_25[39]+inp_26[38];
  assign {FA_cout_551,FA_out_551}=inp_24[42]+inp_25[41]+inp_26[40];
  assign {FA_cout_552,FA_out_552}=inp_24[45]+inp_25[44]+inp_26[43];
  assign {FA_cout_553,FA_out_553}=inp_24[48]+inp_25[47]+inp_26[46];
  assign {FA_cout_554,FA_out_554}=inp_24[51]+inp_25[50]+inp_26[49];
  assign {FA_cout_555,FA_out_555}=inp_24[54]+inp_25[53]+inp_26[52];
  assign {FA_cout_556,FA_out_556}=inp_24[57]+inp_25[56]+inp_26[55];
  assign {FA_cout_557,FA_out_557}=inp_24[60]+inp_25[59]+inp_26[58];
  assign {FA_cout_558,FA_out_558}=inp_24[63]+inp_25[62]+inp_26[61];
  assign {FA_cout_559,FA_out_559}=inp_25[42]+inp_26[41]+inp_27[40];
  assign {FA_cout_560,FA_out_560}=inp_25[45]+inp_26[44]+inp_27[43];
  assign {FA_cout_561,FA_out_561}=inp_25[48]+inp_26[47]+inp_27[46];
  assign {FA_cout_562,FA_out_562}=inp_25[51]+inp_26[50]+inp_27[49];
  assign {FA_cout_563,FA_out_563}=inp_25[54]+inp_26[53]+inp_27[52];
  assign {FA_cout_564,FA_out_564}=inp_25[57]+inp_26[56]+inp_27[55];
  assign {FA_cout_565,FA_out_565}=inp_25[60]+inp_26[59]+inp_27[58];
  assign {FA_cout_566,FA_out_566}=inp_25[63]+inp_26[62]+inp_27[61];
  assign {FA_cout_567,FA_out_567}=inp_26[39]+inp_27[38]+inp_28[37];
  assign {FA_cout_568,FA_out_568}=inp_26[42]+inp_27[41]+inp_28[40];
  assign {FA_cout_569,FA_out_569}=inp_26[45]+inp_27[44]+inp_28[43];
  assign {FA_cout_570,FA_out_570}=inp_26[48]+inp_27[47]+inp_28[46];
  assign {FA_cout_571,FA_out_571}=inp_26[51]+inp_27[50]+inp_28[49];
  assign {FA_cout_572,FA_out_572}=inp_26[54]+inp_27[53]+inp_28[52];
  assign {FA_cout_573,FA_out_573}=inp_26[57]+inp_27[56]+inp_28[55];
  assign {FA_cout_574,FA_out_574}=inp_26[60]+inp_27[59]+inp_28[58];
  assign {FA_cout_575,FA_out_575}=inp_26[63]+inp_27[62]+inp_28[61];
  assign {FA_cout_576,FA_out_576}=inp_27[2]+inp_28[1]+inp_29[0];
  assign {FA_cout_577,FA_out_577}=inp_27[3]+inp_28[2]+inp_29[1];
  assign {FA_cout_578,FA_out_578}=inp_27[4]+inp_28[3]+inp_29[2];
  assign {FA_cout_579,FA_out_579}=inp_27[5]+inp_28[4]+inp_29[3];
  assign {FA_cout_580,FA_out_580}=inp_27[6]+inp_28[5]+inp_29[4];
  assign {FA_cout_581,FA_out_581}=inp_27[7]+inp_28[6]+inp_29[5];
  assign {FA_cout_582,FA_out_582}=inp_27[8]+inp_28[7]+inp_29[6];
  assign {FA_cout_583,FA_out_583}=inp_27[9]+inp_28[8]+inp_29[7];
  assign {FA_cout_584,FA_out_584}=inp_27[10]+inp_28[9]+inp_29[8];
  assign {FA_cout_585,FA_out_585}=inp_27[11]+inp_28[10]+inp_29[9];
  assign {FA_cout_586,FA_out_586}=inp_27[12]+inp_28[11]+inp_29[10];
  assign {FA_cout_587,FA_out_587}=inp_27[13]+inp_28[12]+inp_29[11];
  assign {FA_cout_588,FA_out_588}=inp_27[14]+inp_28[13]+inp_29[12];
  assign {FA_cout_589,FA_out_589}=inp_27[15]+inp_28[14]+inp_29[13];
  assign {FA_cout_590,FA_out_590}=inp_27[16]+inp_28[15]+inp_29[14];
  assign {FA_cout_591,FA_out_591}=inp_27[17]+inp_28[16]+inp_29[15];
  assign {FA_cout_592,FA_out_592}=inp_27[18]+inp_28[17]+inp_29[16];
  assign {FA_cout_593,FA_out_593}=inp_27[19]+inp_28[18]+inp_29[17];
  assign {FA_cout_594,FA_out_594}=inp_27[20]+inp_28[19]+inp_29[18];
  assign {FA_cout_595,FA_out_595}=inp_27[21]+inp_28[20]+inp_29[19];
  assign {FA_cout_596,FA_out_596}=inp_27[22]+inp_28[21]+inp_29[20];
  assign {FA_cout_597,FA_out_597}=inp_27[23]+inp_28[22]+inp_29[21];
  assign {FA_cout_598,FA_out_598}=inp_27[24]+inp_28[23]+inp_29[22];
  assign {FA_cout_599,FA_out_599}=inp_27[25]+inp_28[24]+inp_29[23];
  assign {FA_cout_600,FA_out_600}=inp_27[26]+inp_28[25]+inp_29[24];
  assign {FA_cout_601,FA_out_601}=inp_27[27]+inp_28[26]+inp_29[25];
  assign {FA_cout_602,FA_out_602}=inp_27[28]+inp_28[27]+inp_29[26];
  assign {FA_cout_603,FA_out_603}=inp_27[29]+inp_28[28]+inp_29[27];
  assign {FA_cout_604,FA_out_604}=inp_27[30]+inp_28[29]+inp_29[28];
  assign {FA_cout_605,FA_out_605}=inp_27[31]+inp_28[30]+inp_29[29];
  assign {FA_cout_606,FA_out_606}=inp_27[32]+inp_28[31]+inp_29[30];
  assign {FA_cout_607,FA_out_607}=inp_27[33]+inp_28[32]+inp_29[31];
  assign {FA_cout_608,FA_out_608}=inp_27[34]+inp_28[33]+inp_29[32];
  assign {FA_cout_609,FA_out_609}=inp_27[35]+inp_28[34]+inp_29[33];
  assign {FA_cout_610,FA_out_610}=inp_27[36]+inp_28[35]+inp_29[34];
  assign {FA_cout_611,FA_out_611}=inp_27[37]+inp_28[36]+inp_29[35];
  assign {FA_cout_612,FA_out_612}=inp_27[39]+inp_28[38]+inp_29[37];
  assign {FA_cout_613,FA_out_613}=inp_27[42]+inp_28[41]+inp_29[40];
  assign {FA_cout_614,FA_out_614}=inp_27[45]+inp_28[44]+inp_29[43];
  assign {FA_cout_615,FA_out_615}=inp_27[48]+inp_28[47]+inp_29[46];
  assign {FA_cout_616,FA_out_616}=inp_27[51]+inp_28[50]+inp_29[49];
  assign {FA_cout_617,FA_out_617}=inp_27[54]+inp_28[53]+inp_29[52];
  assign {FA_cout_618,FA_out_618}=inp_27[57]+inp_28[56]+inp_29[55];
  assign {FA_cout_619,FA_out_619}=inp_27[60]+inp_28[59]+inp_29[58];
  assign {FA_cout_620,FA_out_620}=inp_27[63]+inp_28[62]+inp_29[61];
  assign {FA_cout_621,FA_out_621}=inp_28[39]+inp_29[38]+inp_30[37];
  assign {FA_cout_622,FA_out_622}=inp_28[42]+inp_29[41]+inp_30[40];
  assign {FA_cout_623,FA_out_623}=inp_28[45]+inp_29[44]+inp_30[43];
  assign {FA_cout_624,FA_out_624}=inp_28[48]+inp_29[47]+inp_30[46];
  assign {FA_cout_625,FA_out_625}=inp_28[51]+inp_29[50]+inp_30[49];
  assign {FA_cout_626,FA_out_626}=inp_28[54]+inp_29[53]+inp_30[52];
  assign {FA_cout_627,FA_out_627}=inp_28[57]+inp_29[56]+inp_30[55];
  assign {FA_cout_628,FA_out_628}=inp_28[60]+inp_29[59]+inp_30[58];
  assign {FA_cout_629,FA_out_629}=inp_28[63]+inp_29[62]+inp_30[61];
  assign {FA_cout_630,FA_out_630}=inp_29[36]+inp_30[35]+inp_31[34];
  assign {FA_cout_631,FA_out_631}=inp_29[39]+inp_30[38]+inp_31[37];
  assign {FA_cout_632,FA_out_632}=inp_29[42]+inp_30[41]+inp_31[40];
  assign {FA_cout_633,FA_out_633}=inp_29[45]+inp_30[44]+inp_31[43];
  assign {FA_cout_634,FA_out_634}=inp_29[48]+inp_30[47]+inp_31[46];
  assign {FA_cout_635,FA_out_635}=inp_29[51]+inp_30[50]+inp_31[49];
  assign {FA_cout_636,FA_out_636}=inp_29[54]+inp_30[53]+inp_31[52];
  assign {FA_cout_637,FA_out_637}=inp_29[57]+inp_30[56]+inp_31[55];
  assign {FA_cout_638,FA_out_638}=inp_29[60]+inp_30[59]+inp_31[58];
  assign {FA_cout_639,FA_out_639}=inp_29[63]+inp_30[62]+inp_31[61];
  assign {FA_cout_640,FA_out_640}=inp_30[2]+inp_31[1]+inp_32[0];
  assign {FA_cout_641,FA_out_641}=inp_30[3]+inp_31[2]+inp_32[1];
  assign {FA_cout_642,FA_out_642}=inp_30[4]+inp_31[3]+inp_32[2];
  assign {FA_cout_643,FA_out_643}=inp_30[5]+inp_31[4]+inp_32[3];
  assign {FA_cout_644,FA_out_644}=inp_30[6]+inp_31[5]+inp_32[4];
  assign {FA_cout_645,FA_out_645}=inp_30[7]+inp_31[6]+inp_32[5];
  assign {FA_cout_646,FA_out_646}=inp_30[8]+inp_31[7]+inp_32[6];
  assign {FA_cout_647,FA_out_647}=inp_30[9]+inp_31[8]+inp_32[7];
  assign {FA_cout_648,FA_out_648}=inp_30[10]+inp_31[9]+inp_32[8];
  assign {FA_cout_649,FA_out_649}=inp_30[11]+inp_31[10]+inp_32[9];
  assign {FA_cout_650,FA_out_650}=inp_30[12]+inp_31[11]+inp_32[10];
  assign {FA_cout_651,FA_out_651}=inp_30[13]+inp_31[12]+inp_32[11];
  assign {FA_cout_652,FA_out_652}=inp_30[14]+inp_31[13]+inp_32[12];
  assign {FA_cout_653,FA_out_653}=inp_30[15]+inp_31[14]+inp_32[13];
  assign {FA_cout_654,FA_out_654}=inp_30[16]+inp_31[15]+inp_32[14];
  assign {FA_cout_655,FA_out_655}=inp_30[17]+inp_31[16]+inp_32[15];
  assign {FA_cout_656,FA_out_656}=inp_30[18]+inp_31[17]+inp_32[16];
  assign {FA_cout_657,FA_out_657}=inp_30[19]+inp_31[18]+inp_32[17];
  assign {FA_cout_658,FA_out_658}=inp_30[20]+inp_31[19]+inp_32[18];
  assign {FA_cout_659,FA_out_659}=inp_30[21]+inp_31[20]+inp_32[19];
  assign {FA_cout_660,FA_out_660}=inp_30[22]+inp_31[21]+inp_32[20];
  assign {FA_cout_661,FA_out_661}=inp_30[23]+inp_31[22]+inp_32[21];
  assign {FA_cout_662,FA_out_662}=inp_30[24]+inp_31[23]+inp_32[22];
  assign {FA_cout_663,FA_out_663}=inp_30[25]+inp_31[24]+inp_32[23];
  assign {FA_cout_664,FA_out_664}=inp_30[26]+inp_31[25]+inp_32[24];
  assign {FA_cout_665,FA_out_665}=inp_30[27]+inp_31[26]+inp_32[25];
  assign {FA_cout_666,FA_out_666}=inp_30[28]+inp_31[27]+inp_32[26];
  assign {FA_cout_667,FA_out_667}=inp_30[29]+inp_31[28]+inp_32[27];
  assign {FA_cout_668,FA_out_668}=inp_30[30]+inp_31[29]+inp_32[28];
  assign {FA_cout_669,FA_out_669}=inp_30[31]+inp_31[30]+inp_32[29];
  assign {FA_cout_670,FA_out_670}=inp_30[32]+inp_31[31]+inp_32[30];
  assign {FA_cout_671,FA_out_671}=inp_30[33]+inp_31[32]+inp_32[31];
  assign {FA_cout_672,FA_out_672}=inp_30[34]+inp_31[33]+inp_32[32];
  assign {FA_cout_673,FA_out_673}=inp_30[36]+inp_31[35]+inp_32[34];
  assign {FA_cout_674,FA_out_674}=inp_30[39]+inp_31[38]+inp_32[37];
  assign {FA_cout_675,FA_out_675}=inp_30[42]+inp_31[41]+inp_32[40];
  assign {FA_cout_676,FA_out_676}=inp_30[45]+inp_31[44]+inp_32[43];
  assign {FA_cout_677,FA_out_677}=inp_30[48]+inp_31[47]+inp_32[46];
  assign {FA_cout_678,FA_out_678}=inp_30[51]+inp_31[50]+inp_32[49];
  assign {FA_cout_679,FA_out_679}=inp_30[54]+inp_31[53]+inp_32[52];
  assign {FA_cout_680,FA_out_680}=inp_30[57]+inp_31[56]+inp_32[55];
  assign {FA_cout_681,FA_out_681}=inp_30[60]+inp_31[59]+inp_32[58];
  assign {FA_cout_682,FA_out_682}=inp_30[63]+inp_31[62]+inp_32[61];
  assign {FA_cout_683,FA_out_683}=inp_31[36]+inp_32[35]+inp_33[34];
  assign {FA_cout_684,FA_out_684}=inp_31[39]+inp_32[38]+inp_33[37];
  assign {FA_cout_685,FA_out_685}=inp_31[42]+inp_32[41]+inp_33[40];
  assign {FA_cout_686,FA_out_686}=inp_31[45]+inp_32[44]+inp_33[43];
  assign {FA_cout_687,FA_out_687}=inp_31[48]+inp_32[47]+inp_33[46];
  assign {FA_cout_688,FA_out_688}=inp_31[51]+inp_32[50]+inp_33[49];
  assign {FA_cout_689,FA_out_689}=inp_31[54]+inp_32[53]+inp_33[52];
  assign {FA_cout_690,FA_out_690}=inp_31[57]+inp_32[56]+inp_33[55];
  assign {FA_cout_691,FA_out_691}=inp_31[60]+inp_32[59]+inp_33[58];
  assign {FA_cout_692,FA_out_692}=inp_31[63]+inp_32[62]+inp_33[61];
  assign {FA_cout_693,FA_out_693}=inp_32[33]+inp_33[32]+inp_34[31];
  assign {FA_cout_694,FA_out_694}=inp_32[36]+inp_33[35]+inp_34[34];
  assign {FA_cout_695,FA_out_695}=inp_32[39]+inp_33[38]+inp_34[37];
  assign {FA_cout_696,FA_out_696}=inp_32[42]+inp_33[41]+inp_34[40];
  assign {FA_cout_697,FA_out_697}=inp_32[45]+inp_33[44]+inp_34[43];
  assign {FA_cout_698,FA_out_698}=inp_32[48]+inp_33[47]+inp_34[46];
  assign {FA_cout_699,FA_out_699}=inp_32[51]+inp_33[50]+inp_34[49];
  assign {FA_cout_700,FA_out_700}=inp_32[54]+inp_33[53]+inp_34[52];
  assign {FA_cout_701,FA_out_701}=inp_32[57]+inp_33[56]+inp_34[55];
  assign {FA_cout_702,FA_out_702}=inp_32[60]+inp_33[59]+inp_34[58];
  assign {FA_cout_703,FA_out_703}=inp_32[63]+inp_33[62]+inp_34[61];
  assign {FA_cout_704,FA_out_704}=inp_33[2]+inp_34[1]+inp_35[0];
  assign {FA_cout_705,FA_out_705}=inp_33[3]+inp_34[2]+inp_35[1];
  assign {FA_cout_706,FA_out_706}=inp_33[4]+inp_34[3]+inp_35[2];
  assign {FA_cout_707,FA_out_707}=inp_33[5]+inp_34[4]+inp_35[3];
  assign {FA_cout_708,FA_out_708}=inp_33[6]+inp_34[5]+inp_35[4];
  assign {FA_cout_709,FA_out_709}=inp_33[7]+inp_34[6]+inp_35[5];
  assign {FA_cout_710,FA_out_710}=inp_33[8]+inp_34[7]+inp_35[6];
  assign {FA_cout_711,FA_out_711}=inp_33[9]+inp_34[8]+inp_35[7];
  assign {FA_cout_712,FA_out_712}=inp_33[10]+inp_34[9]+inp_35[8];
  assign {FA_cout_713,FA_out_713}=inp_33[11]+inp_34[10]+inp_35[9];
  assign {FA_cout_714,FA_out_714}=inp_33[12]+inp_34[11]+inp_35[10];
  assign {FA_cout_715,FA_out_715}=inp_33[13]+inp_34[12]+inp_35[11];
  assign {FA_cout_716,FA_out_716}=inp_33[14]+inp_34[13]+inp_35[12];
  assign {FA_cout_717,FA_out_717}=inp_33[15]+inp_34[14]+inp_35[13];
  assign {FA_cout_718,FA_out_718}=inp_33[16]+inp_34[15]+inp_35[14];
  assign {FA_cout_719,FA_out_719}=inp_33[17]+inp_34[16]+inp_35[15];
  assign {FA_cout_720,FA_out_720}=inp_33[18]+inp_34[17]+inp_35[16];
  assign {FA_cout_721,FA_out_721}=inp_33[19]+inp_34[18]+inp_35[17];
  assign {FA_cout_722,FA_out_722}=inp_33[20]+inp_34[19]+inp_35[18];
  assign {FA_cout_723,FA_out_723}=inp_33[21]+inp_34[20]+inp_35[19];
  assign {FA_cout_724,FA_out_724}=inp_33[22]+inp_34[21]+inp_35[20];
  assign {FA_cout_725,FA_out_725}=inp_33[23]+inp_34[22]+inp_35[21];
  assign {FA_cout_726,FA_out_726}=inp_33[24]+inp_34[23]+inp_35[22];
  assign {FA_cout_727,FA_out_727}=inp_33[25]+inp_34[24]+inp_35[23];
  assign {FA_cout_728,FA_out_728}=inp_33[26]+inp_34[25]+inp_35[24];
  assign {FA_cout_729,FA_out_729}=inp_33[27]+inp_34[26]+inp_35[25];
  assign {FA_cout_730,FA_out_730}=inp_33[28]+inp_34[27]+inp_35[26];
  assign {FA_cout_731,FA_out_731}=inp_33[29]+inp_34[28]+inp_35[27];
  assign {FA_cout_732,FA_out_732}=inp_33[30]+inp_34[29]+inp_35[28];
  assign {FA_cout_733,FA_out_733}=inp_33[31]+inp_34[30]+inp_35[29];
  assign {FA_cout_734,FA_out_734}=inp_33[33]+inp_34[32]+inp_35[31];
  assign {FA_cout_735,FA_out_735}=inp_33[36]+inp_34[35]+inp_35[34];
  assign {FA_cout_736,FA_out_736}=inp_33[39]+inp_34[38]+inp_35[37];
  assign {FA_cout_737,FA_out_737}=inp_33[42]+inp_34[41]+inp_35[40];
  assign {FA_cout_738,FA_out_738}=inp_33[45]+inp_34[44]+inp_35[43];
  assign {FA_cout_739,FA_out_739}=inp_33[48]+inp_34[47]+inp_35[46];
  assign {FA_cout_740,FA_out_740}=inp_33[51]+inp_34[50]+inp_35[49];
  assign {FA_cout_741,FA_out_741}=inp_33[54]+inp_34[53]+inp_35[52];
  assign {FA_cout_742,FA_out_742}=inp_33[57]+inp_34[56]+inp_35[55];
  assign {FA_cout_743,FA_out_743}=inp_33[60]+inp_34[59]+inp_35[58];
  assign {FA_cout_744,FA_out_744}=inp_33[63]+inp_34[62]+inp_35[61];
  assign {FA_cout_745,FA_out_745}=inp_34[33]+inp_35[32]+inp_36[31];
  assign {FA_cout_746,FA_out_746}=inp_34[36]+inp_35[35]+inp_36[34];
  assign {FA_cout_747,FA_out_747}=inp_34[39]+inp_35[38]+inp_36[37];
  assign {FA_cout_748,FA_out_748}=inp_34[42]+inp_35[41]+inp_36[40];
  assign {FA_cout_749,FA_out_749}=inp_34[45]+inp_35[44]+inp_36[43];
  assign {FA_cout_750,FA_out_750}=inp_34[48]+inp_35[47]+inp_36[46];
  assign {FA_cout_751,FA_out_751}=inp_34[51]+inp_35[50]+inp_36[49];
  assign {FA_cout_752,FA_out_752}=inp_34[54]+inp_35[53]+inp_36[52];
  assign {FA_cout_753,FA_out_753}=inp_34[57]+inp_35[56]+inp_36[55];
  assign {FA_cout_754,FA_out_754}=inp_34[60]+inp_35[59]+inp_36[58];
  assign {FA_cout_755,FA_out_755}=inp_34[63]+inp_35[62]+inp_36[61];
  assign {FA_cout_756,FA_out_756}=inp_35[30]+inp_36[29]+inp_37[28];
  assign {FA_cout_757,FA_out_757}=inp_35[33]+inp_36[32]+inp_37[31];
  assign {FA_cout_758,FA_out_758}=inp_35[36]+inp_36[35]+inp_37[34];
  assign {FA_cout_759,FA_out_759}=inp_35[39]+inp_36[38]+inp_37[37];
  assign {FA_cout_760,FA_out_760}=inp_35[42]+inp_36[41]+inp_37[40];
  assign {FA_cout_761,FA_out_761}=inp_35[45]+inp_36[44]+inp_37[43];
  assign {FA_cout_762,FA_out_762}=inp_35[48]+inp_36[47]+inp_37[46];
  assign {FA_cout_763,FA_out_763}=inp_35[51]+inp_36[50]+inp_37[49];
  assign {FA_cout_764,FA_out_764}=inp_35[54]+inp_36[53]+inp_37[52];
  assign {FA_cout_765,FA_out_765}=inp_35[57]+inp_36[56]+inp_37[55];
  assign {FA_cout_766,FA_out_766}=inp_35[60]+inp_36[59]+inp_37[58];
  assign {FA_cout_767,FA_out_767}=inp_35[63]+inp_36[62]+inp_37[61];
  assign {FA_cout_768,FA_out_768}=inp_36[2]+inp_37[1]+inp_38[0];
  assign {FA_cout_769,FA_out_769}=inp_36[3]+inp_37[2]+inp_38[1];
  assign {FA_cout_770,FA_out_770}=inp_36[4]+inp_37[3]+inp_38[2];
  assign {FA_cout_771,FA_out_771}=inp_36[5]+inp_37[4]+inp_38[3];
  assign {FA_cout_772,FA_out_772}=inp_36[6]+inp_37[5]+inp_38[4];
  assign {FA_cout_773,FA_out_773}=inp_36[7]+inp_37[6]+inp_38[5];
  assign {FA_cout_774,FA_out_774}=inp_36[8]+inp_37[7]+inp_38[6];
  assign {FA_cout_775,FA_out_775}=inp_36[9]+inp_37[8]+inp_38[7];
  assign {FA_cout_776,FA_out_776}=inp_36[10]+inp_37[9]+inp_38[8];
  assign {FA_cout_777,FA_out_777}=inp_36[11]+inp_37[10]+inp_38[9];
  assign {FA_cout_778,FA_out_778}=inp_36[12]+inp_37[11]+inp_38[10];
  assign {FA_cout_779,FA_out_779}=inp_36[13]+inp_37[12]+inp_38[11];
  assign {FA_cout_780,FA_out_780}=inp_36[14]+inp_37[13]+inp_38[12];
  assign {FA_cout_781,FA_out_781}=inp_36[15]+inp_37[14]+inp_38[13];
  assign {FA_cout_782,FA_out_782}=inp_36[16]+inp_37[15]+inp_38[14];
  assign {FA_cout_783,FA_out_783}=inp_36[17]+inp_37[16]+inp_38[15];
  assign {FA_cout_784,FA_out_784}=inp_36[18]+inp_37[17]+inp_38[16];
  assign {FA_cout_785,FA_out_785}=inp_36[19]+inp_37[18]+inp_38[17];
  assign {FA_cout_786,FA_out_786}=inp_36[20]+inp_37[19]+inp_38[18];
  assign {FA_cout_787,FA_out_787}=inp_36[21]+inp_37[20]+inp_38[19];
  assign {FA_cout_788,FA_out_788}=inp_36[22]+inp_37[21]+inp_38[20];
  assign {FA_cout_789,FA_out_789}=inp_36[23]+inp_37[22]+inp_38[21];
  assign {FA_cout_790,FA_out_790}=inp_36[24]+inp_37[23]+inp_38[22];
  assign {FA_cout_791,FA_out_791}=inp_36[25]+inp_37[24]+inp_38[23];
  assign {FA_cout_792,FA_out_792}=inp_36[26]+inp_37[25]+inp_38[24];
  assign {FA_cout_793,FA_out_793}=inp_36[27]+inp_37[26]+inp_38[25];
  assign {FA_cout_794,FA_out_794}=inp_36[28]+inp_37[27]+inp_38[26];
  assign {FA_cout_795,FA_out_795}=inp_36[30]+inp_37[29]+inp_38[28];
  assign {FA_cout_796,FA_out_796}=inp_36[33]+inp_37[32]+inp_38[31];
  assign {FA_cout_797,FA_out_797}=inp_36[36]+inp_37[35]+inp_38[34];
  assign {FA_cout_798,FA_out_798}=inp_36[39]+inp_37[38]+inp_38[37];
  assign {FA_cout_799,FA_out_799}=inp_36[42]+inp_37[41]+inp_38[40];
  assign {FA_cout_800,FA_out_800}=inp_36[45]+inp_37[44]+inp_38[43];
  assign {FA_cout_801,FA_out_801}=inp_36[48]+inp_37[47]+inp_38[46];
  assign {FA_cout_802,FA_out_802}=inp_36[51]+inp_37[50]+inp_38[49];
  assign {FA_cout_803,FA_out_803}=inp_36[54]+inp_37[53]+inp_38[52];
  assign {FA_cout_804,FA_out_804}=inp_36[57]+inp_37[56]+inp_38[55];
  assign {FA_cout_805,FA_out_805}=inp_36[60]+inp_37[59]+inp_38[58];
  assign {FA_cout_806,FA_out_806}=inp_36[63]+inp_37[62]+inp_38[61];
  assign {FA_cout_807,FA_out_807}=inp_37[30]+inp_38[29]+inp_39[28];
  assign {FA_cout_808,FA_out_808}=inp_37[33]+inp_38[32]+inp_39[31];
  assign {FA_cout_809,FA_out_809}=inp_37[36]+inp_38[35]+inp_39[34];
  assign {FA_cout_810,FA_out_810}=inp_37[39]+inp_38[38]+inp_39[37];
  assign {FA_cout_811,FA_out_811}=inp_37[42]+inp_38[41]+inp_39[40];
  assign {FA_cout_812,FA_out_812}=inp_37[45]+inp_38[44]+inp_39[43];
  assign {FA_cout_813,FA_out_813}=inp_37[48]+inp_38[47]+inp_39[46];
  assign {FA_cout_814,FA_out_814}=inp_37[51]+inp_38[50]+inp_39[49];
  assign {FA_cout_815,FA_out_815}=inp_37[54]+inp_38[53]+inp_39[52];
  assign {FA_cout_816,FA_out_816}=inp_37[57]+inp_38[56]+inp_39[55];
  assign {FA_cout_817,FA_out_817}=inp_37[60]+inp_38[59]+inp_39[58];
  assign {FA_cout_818,FA_out_818}=inp_37[63]+inp_38[62]+inp_39[61];
  assign {FA_cout_819,FA_out_819}=inp_38[27]+inp_39[26]+inp_40[25];
  assign {FA_cout_820,FA_out_820}=inp_38[30]+inp_39[29]+inp_40[28];
  assign {FA_cout_821,FA_out_821}=inp_38[33]+inp_39[32]+inp_40[31];
  assign {FA_cout_822,FA_out_822}=inp_38[36]+inp_39[35]+inp_40[34];
  assign {FA_cout_823,FA_out_823}=inp_38[39]+inp_39[38]+inp_40[37];
  assign {FA_cout_824,FA_out_824}=inp_38[42]+inp_39[41]+inp_40[40];
  assign {FA_cout_825,FA_out_825}=inp_38[45]+inp_39[44]+inp_40[43];
  assign {FA_cout_826,FA_out_826}=inp_38[48]+inp_39[47]+inp_40[46];
  assign {FA_cout_827,FA_out_827}=inp_38[51]+inp_39[50]+inp_40[49];
  assign {FA_cout_828,FA_out_828}=inp_38[54]+inp_39[53]+inp_40[52];
  assign {FA_cout_829,FA_out_829}=inp_38[57]+inp_39[56]+inp_40[55];
  assign {FA_cout_830,FA_out_830}=inp_38[60]+inp_39[59]+inp_40[58];
  assign {FA_cout_831,FA_out_831}=inp_38[63]+inp_39[62]+inp_40[61];
  assign {FA_cout_832,FA_out_832}=inp_39[2]+inp_40[1]+inp_41[0];
  assign {FA_cout_833,FA_out_833}=inp_39[3]+inp_40[2]+inp_41[1];
  assign {FA_cout_834,FA_out_834}=inp_39[4]+inp_40[3]+inp_41[2];
  assign {FA_cout_835,FA_out_835}=inp_39[5]+inp_40[4]+inp_41[3];
  assign {FA_cout_836,FA_out_836}=inp_39[6]+inp_40[5]+inp_41[4];
  assign {FA_cout_837,FA_out_837}=inp_39[7]+inp_40[6]+inp_41[5];
  assign {FA_cout_838,FA_out_838}=inp_39[8]+inp_40[7]+inp_41[6];
  assign {FA_cout_839,FA_out_839}=inp_39[9]+inp_40[8]+inp_41[7];
  assign {FA_cout_840,FA_out_840}=inp_39[10]+inp_40[9]+inp_41[8];
  assign {FA_cout_841,FA_out_841}=inp_39[11]+inp_40[10]+inp_41[9];
  assign {FA_cout_842,FA_out_842}=inp_39[12]+inp_40[11]+inp_41[10];
  assign {FA_cout_843,FA_out_843}=inp_39[13]+inp_40[12]+inp_41[11];
  assign {FA_cout_844,FA_out_844}=inp_39[14]+inp_40[13]+inp_41[12];
  assign {FA_cout_845,FA_out_845}=inp_39[15]+inp_40[14]+inp_41[13];
  assign {FA_cout_846,FA_out_846}=inp_39[16]+inp_40[15]+inp_41[14];
  assign {FA_cout_847,FA_out_847}=inp_39[17]+inp_40[16]+inp_41[15];
  assign {FA_cout_848,FA_out_848}=inp_39[18]+inp_40[17]+inp_41[16];
  assign {FA_cout_849,FA_out_849}=inp_39[19]+inp_40[18]+inp_41[17];
  assign {FA_cout_850,FA_out_850}=inp_39[20]+inp_40[19]+inp_41[18];
  assign {FA_cout_851,FA_out_851}=inp_39[21]+inp_40[20]+inp_41[19];
  assign {FA_cout_852,FA_out_852}=inp_39[22]+inp_40[21]+inp_41[20];
  assign {FA_cout_853,FA_out_853}=inp_39[23]+inp_40[22]+inp_41[21];
  assign {FA_cout_854,FA_out_854}=inp_39[24]+inp_40[23]+inp_41[22];
  assign {FA_cout_855,FA_out_855}=inp_39[25]+inp_40[24]+inp_41[23];
  assign {FA_cout_856,FA_out_856}=inp_39[27]+inp_40[26]+inp_41[25];
  assign {FA_cout_857,FA_out_857}=inp_39[30]+inp_40[29]+inp_41[28];
  assign {FA_cout_858,FA_out_858}=inp_39[33]+inp_40[32]+inp_41[31];
  assign {FA_cout_859,FA_out_859}=inp_39[36]+inp_40[35]+inp_41[34];
  assign {FA_cout_860,FA_out_860}=inp_39[39]+inp_40[38]+inp_41[37];
  assign {FA_cout_861,FA_out_861}=inp_39[42]+inp_40[41]+inp_41[40];
  assign {FA_cout_862,FA_out_862}=inp_39[45]+inp_40[44]+inp_41[43];
  assign {FA_cout_863,FA_out_863}=inp_39[48]+inp_40[47]+inp_41[46];
  assign {FA_cout_864,FA_out_864}=inp_39[51]+inp_40[50]+inp_41[49];
  assign {FA_cout_865,FA_out_865}=inp_39[54]+inp_40[53]+inp_41[52];
  assign {FA_cout_866,FA_out_866}=inp_39[57]+inp_40[56]+inp_41[55];
  assign {FA_cout_867,FA_out_867}=inp_39[60]+inp_40[59]+inp_41[58];
  assign {FA_cout_868,FA_out_868}=inp_39[63]+inp_40[62]+inp_41[61];
  assign {FA_cout_869,FA_out_869}=inp_40[27]+inp_41[26]+inp_42[25];
  assign {FA_cout_870,FA_out_870}=inp_40[30]+inp_41[29]+inp_42[28];
  assign {FA_cout_871,FA_out_871}=inp_40[33]+inp_41[32]+inp_42[31];
  assign {FA_cout_872,FA_out_872}=inp_40[36]+inp_41[35]+inp_42[34];
  assign {FA_cout_873,FA_out_873}=inp_40[39]+inp_41[38]+inp_42[37];
  assign {FA_cout_874,FA_out_874}=inp_40[42]+inp_41[41]+inp_42[40];
  assign {FA_cout_875,FA_out_875}=inp_40[45]+inp_41[44]+inp_42[43];
  assign {FA_cout_876,FA_out_876}=inp_40[48]+inp_41[47]+inp_42[46];
  assign {FA_cout_877,FA_out_877}=inp_40[51]+inp_41[50]+inp_42[49];
  assign {FA_cout_878,FA_out_878}=inp_40[54]+inp_41[53]+inp_42[52];
  assign {FA_cout_879,FA_out_879}=inp_40[57]+inp_41[56]+inp_42[55];
  assign {FA_cout_880,FA_out_880}=inp_40[60]+inp_41[59]+inp_42[58];
  assign {FA_cout_881,FA_out_881}=inp_40[63]+inp_41[62]+inp_42[61];
  assign {FA_cout_882,FA_out_882}=inp_41[24]+inp_42[23]+inp_43[22];
  assign {FA_cout_883,FA_out_883}=inp_41[27]+inp_42[26]+inp_43[25];
  assign {FA_cout_884,FA_out_884}=inp_41[30]+inp_42[29]+inp_43[28];
  assign {FA_cout_885,FA_out_885}=inp_41[33]+inp_42[32]+inp_43[31];
  assign {FA_cout_886,FA_out_886}=inp_41[36]+inp_42[35]+inp_43[34];
  assign {FA_cout_887,FA_out_887}=inp_41[39]+inp_42[38]+inp_43[37];
  assign {FA_cout_888,FA_out_888}=inp_41[42]+inp_42[41]+inp_43[40];
  assign {FA_cout_889,FA_out_889}=inp_41[45]+inp_42[44]+inp_43[43];
  assign {FA_cout_890,FA_out_890}=inp_41[48]+inp_42[47]+inp_43[46];
  assign {FA_cout_891,FA_out_891}=inp_41[51]+inp_42[50]+inp_43[49];
  assign {FA_cout_892,FA_out_892}=inp_41[54]+inp_42[53]+inp_43[52];
  assign {FA_cout_893,FA_out_893}=inp_41[57]+inp_42[56]+inp_43[55];
  assign {FA_cout_894,FA_out_894}=inp_41[60]+inp_42[59]+inp_43[58];
  assign {FA_cout_895,FA_out_895}=inp_41[63]+inp_42[62]+inp_43[61];
  assign {FA_cout_896,FA_out_896}=inp_42[2]+inp_43[1]+inp_44[0];
  assign {FA_cout_897,FA_out_897}=inp_42[3]+inp_43[2]+inp_44[1];
  assign {FA_cout_898,FA_out_898}=inp_42[4]+inp_43[3]+inp_44[2];
  assign {FA_cout_899,FA_out_899}=inp_42[5]+inp_43[4]+inp_44[3];
  assign {FA_cout_900,FA_out_900}=inp_42[6]+inp_43[5]+inp_44[4];
  assign {FA_cout_901,FA_out_901}=inp_42[7]+inp_43[6]+inp_44[5];
  assign {FA_cout_902,FA_out_902}=inp_42[8]+inp_43[7]+inp_44[6];
  assign {FA_cout_903,FA_out_903}=inp_42[9]+inp_43[8]+inp_44[7];
  assign {FA_cout_904,FA_out_904}=inp_42[10]+inp_43[9]+inp_44[8];
  assign {FA_cout_905,FA_out_905}=inp_42[11]+inp_43[10]+inp_44[9];
  assign {FA_cout_906,FA_out_906}=inp_42[12]+inp_43[11]+inp_44[10];
  assign {FA_cout_907,FA_out_907}=inp_42[13]+inp_43[12]+inp_44[11];
  assign {FA_cout_908,FA_out_908}=inp_42[14]+inp_43[13]+inp_44[12];
  assign {FA_cout_909,FA_out_909}=inp_42[15]+inp_43[14]+inp_44[13];
  assign {FA_cout_910,FA_out_910}=inp_42[16]+inp_43[15]+inp_44[14];
  assign {FA_cout_911,FA_out_911}=inp_42[17]+inp_43[16]+inp_44[15];
  assign {FA_cout_912,FA_out_912}=inp_42[18]+inp_43[17]+inp_44[16];
  assign {FA_cout_913,FA_out_913}=inp_42[19]+inp_43[18]+inp_44[17];
  assign {FA_cout_914,FA_out_914}=inp_42[20]+inp_43[19]+inp_44[18];
  assign {FA_cout_915,FA_out_915}=inp_42[21]+inp_43[20]+inp_44[19];
  assign {FA_cout_916,FA_out_916}=inp_42[22]+inp_43[21]+inp_44[20];
  assign {FA_cout_917,FA_out_917}=inp_42[24]+inp_43[23]+inp_44[22];
  assign {FA_cout_918,FA_out_918}=inp_42[27]+inp_43[26]+inp_44[25];
  assign {FA_cout_919,FA_out_919}=inp_42[30]+inp_43[29]+inp_44[28];
  assign {FA_cout_920,FA_out_920}=inp_42[33]+inp_43[32]+inp_44[31];
  assign {FA_cout_921,FA_out_921}=inp_42[36]+inp_43[35]+inp_44[34];
  assign {FA_cout_922,FA_out_922}=inp_42[39]+inp_43[38]+inp_44[37];
  assign {FA_cout_923,FA_out_923}=inp_42[42]+inp_43[41]+inp_44[40];
  assign {FA_cout_924,FA_out_924}=inp_42[45]+inp_43[44]+inp_44[43];
  assign {FA_cout_925,FA_out_925}=inp_42[48]+inp_43[47]+inp_44[46];
  assign {FA_cout_926,FA_out_926}=inp_42[51]+inp_43[50]+inp_44[49];
  assign {FA_cout_927,FA_out_927}=inp_42[54]+inp_43[53]+inp_44[52];
  assign {FA_cout_928,FA_out_928}=inp_42[57]+inp_43[56]+inp_44[55];
  assign {FA_cout_929,FA_out_929}=inp_42[60]+inp_43[59]+inp_44[58];
  assign {FA_cout_930,FA_out_930}=inp_42[63]+inp_43[62]+inp_44[61];
  assign {FA_cout_931,FA_out_931}=inp_43[24]+inp_44[23]+inp_45[22];
  assign {FA_cout_932,FA_out_932}=inp_43[27]+inp_44[26]+inp_45[25];
  assign {FA_cout_933,FA_out_933}=inp_43[30]+inp_44[29]+inp_45[28];
  assign {FA_cout_934,FA_out_934}=inp_43[33]+inp_44[32]+inp_45[31];
  assign {FA_cout_935,FA_out_935}=inp_43[36]+inp_44[35]+inp_45[34];
  assign {FA_cout_936,FA_out_936}=inp_43[39]+inp_44[38]+inp_45[37];
  assign {FA_cout_937,FA_out_937}=inp_43[42]+inp_44[41]+inp_45[40];
  assign {FA_cout_938,FA_out_938}=inp_43[45]+inp_44[44]+inp_45[43];
  assign {FA_cout_939,FA_out_939}=inp_43[48]+inp_44[47]+inp_45[46];
  assign {FA_cout_940,FA_out_940}=inp_43[51]+inp_44[50]+inp_45[49];
  assign {FA_cout_941,FA_out_941}=inp_43[54]+inp_44[53]+inp_45[52];
  assign {FA_cout_942,FA_out_942}=inp_43[57]+inp_44[56]+inp_45[55];
  assign {FA_cout_943,FA_out_943}=inp_43[60]+inp_44[59]+inp_45[58];
  assign {FA_cout_944,FA_out_944}=inp_43[63]+inp_44[62]+inp_45[61];
  assign {FA_cout_945,FA_out_945}=inp_44[21]+inp_45[20]+inp_46[19];
  assign {FA_cout_946,FA_out_946}=inp_44[24]+inp_45[23]+inp_46[22];
  assign {FA_cout_947,FA_out_947}=inp_44[27]+inp_45[26]+inp_46[25];
  assign {FA_cout_948,FA_out_948}=inp_44[30]+inp_45[29]+inp_46[28];
  assign {FA_cout_949,FA_out_949}=inp_44[33]+inp_45[32]+inp_46[31];
  assign {FA_cout_950,FA_out_950}=inp_44[36]+inp_45[35]+inp_46[34];
  assign {FA_cout_951,FA_out_951}=inp_44[39]+inp_45[38]+inp_46[37];
  assign {FA_cout_952,FA_out_952}=inp_44[42]+inp_45[41]+inp_46[40];
  assign {FA_cout_953,FA_out_953}=inp_44[45]+inp_45[44]+inp_46[43];
  assign {FA_cout_954,FA_out_954}=inp_44[48]+inp_45[47]+inp_46[46];
  assign {FA_cout_955,FA_out_955}=inp_44[51]+inp_45[50]+inp_46[49];
  assign {FA_cout_956,FA_out_956}=inp_44[54]+inp_45[53]+inp_46[52];
  assign {FA_cout_957,FA_out_957}=inp_44[57]+inp_45[56]+inp_46[55];
  assign {FA_cout_958,FA_out_958}=inp_44[60]+inp_45[59]+inp_46[58];
  assign {FA_cout_959,FA_out_959}=inp_44[63]+inp_45[62]+inp_46[61];
  assign {FA_cout_960,FA_out_960}=inp_45[2]+inp_46[1]+inp_47[0];
  assign {FA_cout_961,FA_out_961}=inp_45[3]+inp_46[2]+inp_47[1];
  assign {FA_cout_962,FA_out_962}=inp_45[4]+inp_46[3]+inp_47[2];
  assign {FA_cout_963,FA_out_963}=inp_45[5]+inp_46[4]+inp_47[3];
  assign {FA_cout_964,FA_out_964}=inp_45[6]+inp_46[5]+inp_47[4];
  assign {FA_cout_965,FA_out_965}=inp_45[7]+inp_46[6]+inp_47[5];
  assign {FA_cout_966,FA_out_966}=inp_45[8]+inp_46[7]+inp_47[6];
  assign {FA_cout_967,FA_out_967}=inp_45[9]+inp_46[8]+inp_47[7];
  assign {FA_cout_968,FA_out_968}=inp_45[10]+inp_46[9]+inp_47[8];
  assign {FA_cout_969,FA_out_969}=inp_45[11]+inp_46[10]+inp_47[9];
  assign {FA_cout_970,FA_out_970}=inp_45[12]+inp_46[11]+inp_47[10];
  assign {FA_cout_971,FA_out_971}=inp_45[13]+inp_46[12]+inp_47[11];
  assign {FA_cout_972,FA_out_972}=inp_45[14]+inp_46[13]+inp_47[12];
  assign {FA_cout_973,FA_out_973}=inp_45[15]+inp_46[14]+inp_47[13];
  assign {FA_cout_974,FA_out_974}=inp_45[16]+inp_46[15]+inp_47[14];
  assign {FA_cout_975,FA_out_975}=inp_45[17]+inp_46[16]+inp_47[15];
  assign {FA_cout_976,FA_out_976}=inp_45[18]+inp_46[17]+inp_47[16];
  assign {FA_cout_977,FA_out_977}=inp_45[19]+inp_46[18]+inp_47[17];
  assign {FA_cout_978,FA_out_978}=inp_45[21]+inp_46[20]+inp_47[19];
  assign {FA_cout_979,FA_out_979}=inp_45[24]+inp_46[23]+inp_47[22];
  assign {FA_cout_980,FA_out_980}=inp_45[27]+inp_46[26]+inp_47[25];
  assign {FA_cout_981,FA_out_981}=inp_45[30]+inp_46[29]+inp_47[28];
  assign {FA_cout_982,FA_out_982}=inp_45[33]+inp_46[32]+inp_47[31];
  assign {FA_cout_983,FA_out_983}=inp_45[36]+inp_46[35]+inp_47[34];
  assign {FA_cout_984,FA_out_984}=inp_45[39]+inp_46[38]+inp_47[37];
  assign {FA_cout_985,FA_out_985}=inp_45[42]+inp_46[41]+inp_47[40];
  assign {FA_cout_986,FA_out_986}=inp_45[45]+inp_46[44]+inp_47[43];
  assign {FA_cout_987,FA_out_987}=inp_45[48]+inp_46[47]+inp_47[46];
  assign {FA_cout_988,FA_out_988}=inp_45[51]+inp_46[50]+inp_47[49];
  assign {FA_cout_989,FA_out_989}=inp_45[54]+inp_46[53]+inp_47[52];
  assign {FA_cout_990,FA_out_990}=inp_45[57]+inp_46[56]+inp_47[55];
  assign {FA_cout_991,FA_out_991}=inp_45[60]+inp_46[59]+inp_47[58];
  assign {FA_cout_992,FA_out_992}=inp_45[63]+inp_46[62]+inp_47[61];
  assign {FA_cout_993,FA_out_993}=inp_46[21]+inp_47[20]+inp_48[19];
  assign {FA_cout_994,FA_out_994}=inp_46[24]+inp_47[23]+inp_48[22];
  assign {FA_cout_995,FA_out_995}=inp_46[27]+inp_47[26]+inp_48[25];
  assign {FA_cout_996,FA_out_996}=inp_46[30]+inp_47[29]+inp_48[28];
  assign {FA_cout_997,FA_out_997}=inp_46[33]+inp_47[32]+inp_48[31];
  assign {FA_cout_998,FA_out_998}=inp_46[36]+inp_47[35]+inp_48[34];
  assign {FA_cout_999,FA_out_999}=inp_46[39]+inp_47[38]+inp_48[37];
  assign {FA_cout_1000,FA_out_1000}=inp_46[42]+inp_47[41]+inp_48[40];
  assign {FA_cout_1001,FA_out_1001}=inp_46[45]+inp_47[44]+inp_48[43];
  assign {FA_cout_1002,FA_out_1002}=inp_46[48]+inp_47[47]+inp_48[46];
  assign {FA_cout_1003,FA_out_1003}=inp_46[51]+inp_47[50]+inp_48[49];
  assign {FA_cout_1004,FA_out_1004}=inp_46[54]+inp_47[53]+inp_48[52];
  assign {FA_cout_1005,FA_out_1005}=inp_46[57]+inp_47[56]+inp_48[55];
  assign {FA_cout_1006,FA_out_1006}=inp_46[60]+inp_47[59]+inp_48[58];
  assign {FA_cout_1007,FA_out_1007}=inp_46[63]+inp_47[62]+inp_48[61];
  assign {FA_cout_1008,FA_out_1008}=inp_47[18]+inp_48[17]+inp_49[16];
  assign {FA_cout_1009,FA_out_1009}=inp_47[21]+inp_48[20]+inp_49[19];
  assign {FA_cout_1010,FA_out_1010}=inp_47[24]+inp_48[23]+inp_49[22];
  assign {FA_cout_1011,FA_out_1011}=inp_47[27]+inp_48[26]+inp_49[25];
  assign {FA_cout_1012,FA_out_1012}=inp_47[30]+inp_48[29]+inp_49[28];
  assign {FA_cout_1013,FA_out_1013}=inp_47[33]+inp_48[32]+inp_49[31];
  assign {FA_cout_1014,FA_out_1014}=inp_47[36]+inp_48[35]+inp_49[34];
  assign {FA_cout_1015,FA_out_1015}=inp_47[39]+inp_48[38]+inp_49[37];
  assign {FA_cout_1016,FA_out_1016}=inp_47[42]+inp_48[41]+inp_49[40];
  assign {FA_cout_1017,FA_out_1017}=inp_47[45]+inp_48[44]+inp_49[43];
  assign {FA_cout_1018,FA_out_1018}=inp_47[48]+inp_48[47]+inp_49[46];
  assign {FA_cout_1019,FA_out_1019}=inp_47[51]+inp_48[50]+inp_49[49];
  assign {FA_cout_1020,FA_out_1020}=inp_47[54]+inp_48[53]+inp_49[52];
  assign {FA_cout_1021,FA_out_1021}=inp_47[57]+inp_48[56]+inp_49[55];
  assign {FA_cout_1022,FA_out_1022}=inp_47[60]+inp_48[59]+inp_49[58];
  assign {FA_cout_1023,FA_out_1023}=inp_47[63]+inp_48[62]+inp_49[61];
  assign {FA_cout_1024,FA_out_1024}=inp_48[2]+inp_49[1]+inp_50[0];
  assign {FA_cout_1025,FA_out_1025}=inp_48[3]+inp_49[2]+inp_50[1];
  assign {FA_cout_1026,FA_out_1026}=inp_48[4]+inp_49[3]+inp_50[2];
  assign {FA_cout_1027,FA_out_1027}=inp_48[5]+inp_49[4]+inp_50[3];
  assign {FA_cout_1028,FA_out_1028}=inp_48[6]+inp_49[5]+inp_50[4];
  assign {FA_cout_1029,FA_out_1029}=inp_48[7]+inp_49[6]+inp_50[5];
  assign {FA_cout_1030,FA_out_1030}=inp_48[8]+inp_49[7]+inp_50[6];
  assign {FA_cout_1031,FA_out_1031}=inp_48[9]+inp_49[8]+inp_50[7];
  assign {FA_cout_1032,FA_out_1032}=inp_48[10]+inp_49[9]+inp_50[8];
  assign {FA_cout_1033,FA_out_1033}=inp_48[11]+inp_49[10]+inp_50[9];
  assign {FA_cout_1034,FA_out_1034}=inp_48[12]+inp_49[11]+inp_50[10];
  assign {FA_cout_1035,FA_out_1035}=inp_48[13]+inp_49[12]+inp_50[11];
  assign {FA_cout_1036,FA_out_1036}=inp_48[14]+inp_49[13]+inp_50[12];
  assign {FA_cout_1037,FA_out_1037}=inp_48[15]+inp_49[14]+inp_50[13];
  assign {FA_cout_1038,FA_out_1038}=inp_48[16]+inp_49[15]+inp_50[14];
  assign {FA_cout_1039,FA_out_1039}=inp_48[18]+inp_49[17]+inp_50[16];
  assign {FA_cout_1040,FA_out_1040}=inp_48[21]+inp_49[20]+inp_50[19];
  assign {FA_cout_1041,FA_out_1041}=inp_48[24]+inp_49[23]+inp_50[22];
  assign {FA_cout_1042,FA_out_1042}=inp_48[27]+inp_49[26]+inp_50[25];
  assign {FA_cout_1043,FA_out_1043}=inp_48[30]+inp_49[29]+inp_50[28];
  assign {FA_cout_1044,FA_out_1044}=inp_48[33]+inp_49[32]+inp_50[31];
  assign {FA_cout_1045,FA_out_1045}=inp_48[36]+inp_49[35]+inp_50[34];
  assign {FA_cout_1046,FA_out_1046}=inp_48[39]+inp_49[38]+inp_50[37];
  assign {FA_cout_1047,FA_out_1047}=inp_48[42]+inp_49[41]+inp_50[40];
  assign {FA_cout_1048,FA_out_1048}=inp_48[45]+inp_49[44]+inp_50[43];
  assign {FA_cout_1049,FA_out_1049}=inp_48[48]+inp_49[47]+inp_50[46];
  assign {FA_cout_1050,FA_out_1050}=inp_48[51]+inp_49[50]+inp_50[49];
  assign {FA_cout_1051,FA_out_1051}=inp_48[54]+inp_49[53]+inp_50[52];
  assign {FA_cout_1052,FA_out_1052}=inp_48[57]+inp_49[56]+inp_50[55];
  assign {FA_cout_1053,FA_out_1053}=inp_48[60]+inp_49[59]+inp_50[58];
  assign {FA_cout_1054,FA_out_1054}=inp_48[63]+inp_49[62]+inp_50[61];
  assign {FA_cout_1055,FA_out_1055}=inp_49[18]+inp_50[17]+inp_51[16];
  assign {FA_cout_1056,FA_out_1056}=inp_49[21]+inp_50[20]+inp_51[19];
  assign {FA_cout_1057,FA_out_1057}=inp_49[24]+inp_50[23]+inp_51[22];
  assign {FA_cout_1058,FA_out_1058}=inp_49[27]+inp_50[26]+inp_51[25];
  assign {FA_cout_1059,FA_out_1059}=inp_49[30]+inp_50[29]+inp_51[28];
  assign {FA_cout_1060,FA_out_1060}=inp_49[33]+inp_50[32]+inp_51[31];
  assign {FA_cout_1061,FA_out_1061}=inp_49[36]+inp_50[35]+inp_51[34];
  assign {FA_cout_1062,FA_out_1062}=inp_49[39]+inp_50[38]+inp_51[37];
  assign {FA_cout_1063,FA_out_1063}=inp_49[42]+inp_50[41]+inp_51[40];
  assign {FA_cout_1064,FA_out_1064}=inp_49[45]+inp_50[44]+inp_51[43];
  assign {FA_cout_1065,FA_out_1065}=inp_49[48]+inp_50[47]+inp_51[46];
  assign {FA_cout_1066,FA_out_1066}=inp_49[51]+inp_50[50]+inp_51[49];
  assign {FA_cout_1067,FA_out_1067}=inp_49[54]+inp_50[53]+inp_51[52];
  assign {FA_cout_1068,FA_out_1068}=inp_49[57]+inp_50[56]+inp_51[55];
  assign {FA_cout_1069,FA_out_1069}=inp_49[60]+inp_50[59]+inp_51[58];
  assign {FA_cout_1070,FA_out_1070}=inp_49[63]+inp_50[62]+inp_51[61];
  assign {FA_cout_1071,FA_out_1071}=inp_50[15]+inp_51[14]+inp_52[13];
  assign {FA_cout_1072,FA_out_1072}=inp_50[18]+inp_51[17]+inp_52[16];
  assign {FA_cout_1073,FA_out_1073}=inp_50[21]+inp_51[20]+inp_52[19];
  assign {FA_cout_1074,FA_out_1074}=inp_50[24]+inp_51[23]+inp_52[22];
  assign {FA_cout_1075,FA_out_1075}=inp_50[27]+inp_51[26]+inp_52[25];
  assign {FA_cout_1076,FA_out_1076}=inp_50[30]+inp_51[29]+inp_52[28];
  assign {FA_cout_1077,FA_out_1077}=inp_50[33]+inp_51[32]+inp_52[31];
  assign {FA_cout_1078,FA_out_1078}=inp_50[36]+inp_51[35]+inp_52[34];
  assign {FA_cout_1079,FA_out_1079}=inp_50[39]+inp_51[38]+inp_52[37];
  assign {FA_cout_1080,FA_out_1080}=inp_50[42]+inp_51[41]+inp_52[40];
  assign {FA_cout_1081,FA_out_1081}=inp_50[45]+inp_51[44]+inp_52[43];
  assign {FA_cout_1082,FA_out_1082}=inp_50[48]+inp_51[47]+inp_52[46];
  assign {FA_cout_1083,FA_out_1083}=inp_50[51]+inp_51[50]+inp_52[49];
  assign {FA_cout_1084,FA_out_1084}=inp_50[54]+inp_51[53]+inp_52[52];
  assign {FA_cout_1085,FA_out_1085}=inp_50[57]+inp_51[56]+inp_52[55];
  assign {FA_cout_1086,FA_out_1086}=inp_50[60]+inp_51[59]+inp_52[58];
  assign {FA_cout_1087,FA_out_1087}=inp_50[63]+inp_51[62]+inp_52[61];
  assign {FA_cout_1088,FA_out_1088}=inp_51[2]+inp_52[1]+inp_53[0];
  assign {FA_cout_1089,FA_out_1089}=inp_51[3]+inp_52[2]+inp_53[1];
  assign {FA_cout_1090,FA_out_1090}=inp_51[4]+inp_52[3]+inp_53[2];
  assign {FA_cout_1091,FA_out_1091}=inp_51[5]+inp_52[4]+inp_53[3];
  assign {FA_cout_1092,FA_out_1092}=inp_51[6]+inp_52[5]+inp_53[4];
  assign {FA_cout_1093,FA_out_1093}=inp_51[7]+inp_52[6]+inp_53[5];
  assign {FA_cout_1094,FA_out_1094}=inp_51[8]+inp_52[7]+inp_53[6];
  assign {FA_cout_1095,FA_out_1095}=inp_51[9]+inp_52[8]+inp_53[7];
  assign {FA_cout_1096,FA_out_1096}=inp_51[10]+inp_52[9]+inp_53[8];
  assign {FA_cout_1097,FA_out_1097}=inp_51[11]+inp_52[10]+inp_53[9];
  assign {FA_cout_1098,FA_out_1098}=inp_51[12]+inp_52[11]+inp_53[10];
  assign {FA_cout_1099,FA_out_1099}=inp_51[13]+inp_52[12]+inp_53[11];
  assign {FA_cout_1100,FA_out_1100}=inp_51[15]+inp_52[14]+inp_53[13];
  assign {FA_cout_1101,FA_out_1101}=inp_51[18]+inp_52[17]+inp_53[16];
  assign {FA_cout_1102,FA_out_1102}=inp_51[21]+inp_52[20]+inp_53[19];
  assign {FA_cout_1103,FA_out_1103}=inp_51[24]+inp_52[23]+inp_53[22];
  assign {FA_cout_1104,FA_out_1104}=inp_51[27]+inp_52[26]+inp_53[25];
  assign {FA_cout_1105,FA_out_1105}=inp_51[30]+inp_52[29]+inp_53[28];
  assign {FA_cout_1106,FA_out_1106}=inp_51[33]+inp_52[32]+inp_53[31];
  assign {FA_cout_1107,FA_out_1107}=inp_51[36]+inp_52[35]+inp_53[34];
  assign {FA_cout_1108,FA_out_1108}=inp_51[39]+inp_52[38]+inp_53[37];
  assign {FA_cout_1109,FA_out_1109}=inp_51[42]+inp_52[41]+inp_53[40];
  assign {FA_cout_1110,FA_out_1110}=inp_51[45]+inp_52[44]+inp_53[43];
  assign {FA_cout_1111,FA_out_1111}=inp_51[48]+inp_52[47]+inp_53[46];
  assign {FA_cout_1112,FA_out_1112}=inp_51[51]+inp_52[50]+inp_53[49];
  assign {FA_cout_1113,FA_out_1113}=inp_51[54]+inp_52[53]+inp_53[52];
  assign {FA_cout_1114,FA_out_1114}=inp_51[57]+inp_52[56]+inp_53[55];
  assign {FA_cout_1115,FA_out_1115}=inp_51[60]+inp_52[59]+inp_53[58];
  assign {FA_cout_1116,FA_out_1116}=inp_51[63]+inp_52[62]+inp_53[61];
  assign {FA_cout_1117,FA_out_1117}=inp_52[15]+inp_53[14]+inp_54[13];
  assign {FA_cout_1118,FA_out_1118}=inp_52[18]+inp_53[17]+inp_54[16];
  assign {FA_cout_1119,FA_out_1119}=inp_52[21]+inp_53[20]+inp_54[19];
  assign {FA_cout_1120,FA_out_1120}=inp_52[24]+inp_53[23]+inp_54[22];
  assign {FA_cout_1121,FA_out_1121}=inp_52[27]+inp_53[26]+inp_54[25];
  assign {FA_cout_1122,FA_out_1122}=inp_52[30]+inp_53[29]+inp_54[28];
  assign {FA_cout_1123,FA_out_1123}=inp_52[33]+inp_53[32]+inp_54[31];
  assign {FA_cout_1124,FA_out_1124}=inp_52[36]+inp_53[35]+inp_54[34];
  assign {FA_cout_1125,FA_out_1125}=inp_52[39]+inp_53[38]+inp_54[37];
  assign {FA_cout_1126,FA_out_1126}=inp_52[42]+inp_53[41]+inp_54[40];
  assign {FA_cout_1127,FA_out_1127}=inp_52[45]+inp_53[44]+inp_54[43];
  assign {FA_cout_1128,FA_out_1128}=inp_52[48]+inp_53[47]+inp_54[46];
  assign {FA_cout_1129,FA_out_1129}=inp_52[51]+inp_53[50]+inp_54[49];
  assign {FA_cout_1130,FA_out_1130}=inp_52[54]+inp_53[53]+inp_54[52];
  assign {FA_cout_1131,FA_out_1131}=inp_52[57]+inp_53[56]+inp_54[55];
  assign {FA_cout_1132,FA_out_1132}=inp_52[60]+inp_53[59]+inp_54[58];
  assign {FA_cout_1133,FA_out_1133}=inp_52[63]+inp_53[62]+inp_54[61];
  assign {FA_cout_1134,FA_out_1134}=inp_53[12]+inp_54[11]+inp_55[10];
  assign {FA_cout_1135,FA_out_1135}=inp_53[15]+inp_54[14]+inp_55[13];
  assign {FA_cout_1136,FA_out_1136}=inp_53[18]+inp_54[17]+inp_55[16];
  assign {FA_cout_1137,FA_out_1137}=inp_53[21]+inp_54[20]+inp_55[19];
  assign {FA_cout_1138,FA_out_1138}=inp_53[24]+inp_54[23]+inp_55[22];
  assign {FA_cout_1139,FA_out_1139}=inp_53[27]+inp_54[26]+inp_55[25];
  assign {FA_cout_1140,FA_out_1140}=inp_53[30]+inp_54[29]+inp_55[28];
  assign {FA_cout_1141,FA_out_1141}=inp_53[33]+inp_54[32]+inp_55[31];
  assign {FA_cout_1142,FA_out_1142}=inp_53[36]+inp_54[35]+inp_55[34];
  assign {FA_cout_1143,FA_out_1143}=inp_53[39]+inp_54[38]+inp_55[37];
  assign {FA_cout_1144,FA_out_1144}=inp_53[42]+inp_54[41]+inp_55[40];
  assign {FA_cout_1145,FA_out_1145}=inp_53[45]+inp_54[44]+inp_55[43];
  assign {FA_cout_1146,FA_out_1146}=inp_53[48]+inp_54[47]+inp_55[46];
  assign {FA_cout_1147,FA_out_1147}=inp_53[51]+inp_54[50]+inp_55[49];
  assign {FA_cout_1148,FA_out_1148}=inp_53[54]+inp_54[53]+inp_55[52];
  assign {FA_cout_1149,FA_out_1149}=inp_53[57]+inp_54[56]+inp_55[55];
  assign {FA_cout_1150,FA_out_1150}=inp_53[60]+inp_54[59]+inp_55[58];
  assign {FA_cout_1151,FA_out_1151}=inp_53[63]+inp_54[62]+inp_55[61];
  assign {FA_cout_1152,FA_out_1152}=inp_54[2]+inp_55[1]+inp_56[0];
  assign {FA_cout_1153,FA_out_1153}=inp_54[3]+inp_55[2]+inp_56[1];
  assign {FA_cout_1154,FA_out_1154}=inp_54[4]+inp_55[3]+inp_56[2];
  assign {FA_cout_1155,FA_out_1155}=inp_54[5]+inp_55[4]+inp_56[3];
  assign {FA_cout_1156,FA_out_1156}=inp_54[6]+inp_55[5]+inp_56[4];
  assign {FA_cout_1157,FA_out_1157}=inp_54[7]+inp_55[6]+inp_56[5];
  assign {FA_cout_1158,FA_out_1158}=inp_54[8]+inp_55[7]+inp_56[6];
  assign {FA_cout_1159,FA_out_1159}=inp_54[9]+inp_55[8]+inp_56[7];
  assign {FA_cout_1160,FA_out_1160}=inp_54[10]+inp_55[9]+inp_56[8];
  assign {FA_cout_1161,FA_out_1161}=inp_54[12]+inp_55[11]+inp_56[10];
  assign {FA_cout_1162,FA_out_1162}=inp_54[15]+inp_55[14]+inp_56[13];
  assign {FA_cout_1163,FA_out_1163}=inp_54[18]+inp_55[17]+inp_56[16];
  assign {FA_cout_1164,FA_out_1164}=inp_54[21]+inp_55[20]+inp_56[19];
  assign {FA_cout_1165,FA_out_1165}=inp_54[24]+inp_55[23]+inp_56[22];
  assign {FA_cout_1166,FA_out_1166}=inp_54[27]+inp_55[26]+inp_56[25];
  assign {FA_cout_1167,FA_out_1167}=inp_54[30]+inp_55[29]+inp_56[28];
  assign {FA_cout_1168,FA_out_1168}=inp_54[33]+inp_55[32]+inp_56[31];
  assign {FA_cout_1169,FA_out_1169}=inp_54[36]+inp_55[35]+inp_56[34];
  assign {FA_cout_1170,FA_out_1170}=inp_54[39]+inp_55[38]+inp_56[37];
  assign {FA_cout_1171,FA_out_1171}=inp_54[42]+inp_55[41]+inp_56[40];
  assign {FA_cout_1172,FA_out_1172}=inp_54[45]+inp_55[44]+inp_56[43];
  assign {FA_cout_1173,FA_out_1173}=inp_54[48]+inp_55[47]+inp_56[46];
  assign {FA_cout_1174,FA_out_1174}=inp_54[51]+inp_55[50]+inp_56[49];
  assign {FA_cout_1175,FA_out_1175}=inp_54[54]+inp_55[53]+inp_56[52];
  assign {FA_cout_1176,FA_out_1176}=inp_54[57]+inp_55[56]+inp_56[55];
  assign {FA_cout_1177,FA_out_1177}=inp_54[60]+inp_55[59]+inp_56[58];
  assign {FA_cout_1178,FA_out_1178}=inp_54[63]+inp_55[62]+inp_56[61];
  assign {FA_cout_1179,FA_out_1179}=inp_55[12]+inp_56[11]+inp_57[10];
  assign {FA_cout_1180,FA_out_1180}=inp_55[15]+inp_56[14]+inp_57[13];
  assign {FA_cout_1181,FA_out_1181}=inp_55[18]+inp_56[17]+inp_57[16];
  assign {FA_cout_1182,FA_out_1182}=inp_55[21]+inp_56[20]+inp_57[19];
  assign {FA_cout_1183,FA_out_1183}=inp_55[24]+inp_56[23]+inp_57[22];
  assign {FA_cout_1184,FA_out_1184}=inp_55[27]+inp_56[26]+inp_57[25];
  assign {FA_cout_1185,FA_out_1185}=inp_55[30]+inp_56[29]+inp_57[28];
  assign {FA_cout_1186,FA_out_1186}=inp_55[33]+inp_56[32]+inp_57[31];
  assign {FA_cout_1187,FA_out_1187}=inp_55[36]+inp_56[35]+inp_57[34];
  assign {FA_cout_1188,FA_out_1188}=inp_55[39]+inp_56[38]+inp_57[37];
  assign {FA_cout_1189,FA_out_1189}=inp_55[42]+inp_56[41]+inp_57[40];
  assign {FA_cout_1190,FA_out_1190}=inp_55[45]+inp_56[44]+inp_57[43];
  assign {FA_cout_1191,FA_out_1191}=inp_55[48]+inp_56[47]+inp_57[46];
  assign {FA_cout_1192,FA_out_1192}=inp_55[51]+inp_56[50]+inp_57[49];
  assign {FA_cout_1193,FA_out_1193}=inp_55[54]+inp_56[53]+inp_57[52];
  assign {FA_cout_1194,FA_out_1194}=inp_55[57]+inp_56[56]+inp_57[55];
  assign {FA_cout_1195,FA_out_1195}=inp_55[60]+inp_56[59]+inp_57[58];
  assign {FA_cout_1196,FA_out_1196}=inp_55[63]+inp_56[62]+inp_57[61];
  assign {FA_cout_1197,FA_out_1197}=inp_56[9]+inp_57[8]+inp_58[7];
  assign {FA_cout_1198,FA_out_1198}=inp_56[12]+inp_57[11]+inp_58[10];
  assign {FA_cout_1199,FA_out_1199}=inp_56[15]+inp_57[14]+inp_58[13];
  assign {FA_cout_1200,FA_out_1200}=inp_56[18]+inp_57[17]+inp_58[16];
  assign {FA_cout_1201,FA_out_1201}=inp_56[21]+inp_57[20]+inp_58[19];
  assign {FA_cout_1202,FA_out_1202}=inp_56[24]+inp_57[23]+inp_58[22];
  assign {FA_cout_1203,FA_out_1203}=inp_56[27]+inp_57[26]+inp_58[25];
  assign {FA_cout_1204,FA_out_1204}=inp_56[30]+inp_57[29]+inp_58[28];
  assign {FA_cout_1205,FA_out_1205}=inp_56[33]+inp_57[32]+inp_58[31];
  assign {FA_cout_1206,FA_out_1206}=inp_56[36]+inp_57[35]+inp_58[34];
  assign {FA_cout_1207,FA_out_1207}=inp_56[39]+inp_57[38]+inp_58[37];
  assign {FA_cout_1208,FA_out_1208}=inp_56[42]+inp_57[41]+inp_58[40];
  assign {FA_cout_1209,FA_out_1209}=inp_56[45]+inp_57[44]+inp_58[43];
  assign {FA_cout_1210,FA_out_1210}=inp_56[48]+inp_57[47]+inp_58[46];
  assign {FA_cout_1211,FA_out_1211}=inp_56[51]+inp_57[50]+inp_58[49];
  assign {FA_cout_1212,FA_out_1212}=inp_56[54]+inp_57[53]+inp_58[52];
  assign {FA_cout_1213,FA_out_1213}=inp_56[57]+inp_57[56]+inp_58[55];
  assign {FA_cout_1214,FA_out_1214}=inp_56[60]+inp_57[59]+inp_58[58];
  assign {FA_cout_1215,FA_out_1215}=inp_56[63]+inp_57[62]+inp_58[61];
  assign {FA_cout_1216,FA_out_1216}=inp_57[2]+inp_58[1]+inp_59[0];
  assign {FA_cout_1217,FA_out_1217}=inp_57[3]+inp_58[2]+inp_59[1];
  assign {FA_cout_1218,FA_out_1218}=inp_57[4]+inp_58[3]+inp_59[2];
  assign {FA_cout_1219,FA_out_1219}=inp_57[5]+inp_58[4]+inp_59[3];
  assign {FA_cout_1220,FA_out_1220}=inp_57[6]+inp_58[5]+inp_59[4];
  assign {FA_cout_1221,FA_out_1221}=inp_57[7]+inp_58[6]+inp_59[5];
  assign {FA_cout_1222,FA_out_1222}=inp_57[9]+inp_58[8]+inp_59[7];
  assign {FA_cout_1223,FA_out_1223}=inp_57[12]+inp_58[11]+inp_59[10];
  assign {FA_cout_1224,FA_out_1224}=inp_57[15]+inp_58[14]+inp_59[13];
  assign {FA_cout_1225,FA_out_1225}=inp_57[18]+inp_58[17]+inp_59[16];
  assign {FA_cout_1226,FA_out_1226}=inp_57[21]+inp_58[20]+inp_59[19];
  assign {FA_cout_1227,FA_out_1227}=inp_57[24]+inp_58[23]+inp_59[22];
  assign {FA_cout_1228,FA_out_1228}=inp_57[27]+inp_58[26]+inp_59[25];
  assign {FA_cout_1229,FA_out_1229}=inp_57[30]+inp_58[29]+inp_59[28];
  assign {FA_cout_1230,FA_out_1230}=inp_57[33]+inp_58[32]+inp_59[31];
  assign {FA_cout_1231,FA_out_1231}=inp_57[36]+inp_58[35]+inp_59[34];
  assign {FA_cout_1232,FA_out_1232}=inp_57[39]+inp_58[38]+inp_59[37];
  assign {FA_cout_1233,FA_out_1233}=inp_57[42]+inp_58[41]+inp_59[40];
  assign {FA_cout_1234,FA_out_1234}=inp_57[45]+inp_58[44]+inp_59[43];
  assign {FA_cout_1235,FA_out_1235}=inp_57[48]+inp_58[47]+inp_59[46];
  assign {FA_cout_1236,FA_out_1236}=inp_57[51]+inp_58[50]+inp_59[49];
  assign {FA_cout_1237,FA_out_1237}=inp_57[54]+inp_58[53]+inp_59[52];
  assign {FA_cout_1238,FA_out_1238}=inp_57[57]+inp_58[56]+inp_59[55];
  assign {FA_cout_1239,FA_out_1239}=inp_57[60]+inp_58[59]+inp_59[58];
  assign {FA_cout_1240,FA_out_1240}=inp_57[63]+inp_58[62]+inp_59[61];
  assign {FA_cout_1241,FA_out_1241}=inp_58[9]+inp_59[8]+inp_60[7];
  assign {FA_cout_1242,FA_out_1242}=inp_58[12]+inp_59[11]+inp_60[10];
  assign {FA_cout_1243,FA_out_1243}=inp_58[15]+inp_59[14]+inp_60[13];
  assign {FA_cout_1244,FA_out_1244}=inp_58[18]+inp_59[17]+inp_60[16];
  assign {FA_cout_1245,FA_out_1245}=inp_58[21]+inp_59[20]+inp_60[19];
  assign {FA_cout_1246,FA_out_1246}=inp_58[24]+inp_59[23]+inp_60[22];
  assign {FA_cout_1247,FA_out_1247}=inp_58[27]+inp_59[26]+inp_60[25];
  assign {FA_cout_1248,FA_out_1248}=inp_58[30]+inp_59[29]+inp_60[28];
  assign {FA_cout_1249,FA_out_1249}=inp_58[33]+inp_59[32]+inp_60[31];
  assign {FA_cout_1250,FA_out_1250}=inp_58[36]+inp_59[35]+inp_60[34];
  assign {FA_cout_1251,FA_out_1251}=inp_58[39]+inp_59[38]+inp_60[37];
  assign {FA_cout_1252,FA_out_1252}=inp_58[42]+inp_59[41]+inp_60[40];
  assign {FA_cout_1253,FA_out_1253}=inp_58[45]+inp_59[44]+inp_60[43];
  assign {FA_cout_1254,FA_out_1254}=inp_58[48]+inp_59[47]+inp_60[46];
  assign {FA_cout_1255,FA_out_1255}=inp_58[51]+inp_59[50]+inp_60[49];
  assign {FA_cout_1256,FA_out_1256}=inp_58[54]+inp_59[53]+inp_60[52];
  assign {FA_cout_1257,FA_out_1257}=inp_58[57]+inp_59[56]+inp_60[55];
  assign {FA_cout_1258,FA_out_1258}=inp_58[60]+inp_59[59]+inp_60[58];
  assign {FA_cout_1259,FA_out_1259}=inp_58[63]+inp_59[62]+inp_60[61];
  assign {FA_cout_1260,FA_out_1260}=inp_59[6]+inp_60[5]+inp_61[4];
  assign {FA_cout_1261,FA_out_1261}=inp_59[9]+inp_60[8]+inp_61[7];
  assign {FA_cout_1262,FA_out_1262}=inp_59[12]+inp_60[11]+inp_61[10];
  assign {FA_cout_1263,FA_out_1263}=inp_59[15]+inp_60[14]+inp_61[13];
  assign {FA_cout_1264,FA_out_1264}=inp_59[18]+inp_60[17]+inp_61[16];
  assign {FA_cout_1265,FA_out_1265}=inp_59[21]+inp_60[20]+inp_61[19];
  assign {FA_cout_1266,FA_out_1266}=inp_59[24]+inp_60[23]+inp_61[22];
  assign {FA_cout_1267,FA_out_1267}=inp_59[27]+inp_60[26]+inp_61[25];
  assign {FA_cout_1268,FA_out_1268}=inp_59[30]+inp_60[29]+inp_61[28];
  assign {FA_cout_1269,FA_out_1269}=inp_59[33]+inp_60[32]+inp_61[31];
  assign {FA_cout_1270,FA_out_1270}=inp_59[36]+inp_60[35]+inp_61[34];
  assign {FA_cout_1271,FA_out_1271}=inp_59[39]+inp_60[38]+inp_61[37];
  assign {FA_cout_1272,FA_out_1272}=inp_59[42]+inp_60[41]+inp_61[40];
  assign {FA_cout_1273,FA_out_1273}=inp_59[45]+inp_60[44]+inp_61[43];
  assign {FA_cout_1274,FA_out_1274}=inp_59[48]+inp_60[47]+inp_61[46];
  assign {FA_cout_1275,FA_out_1275}=inp_59[51]+inp_60[50]+inp_61[49];
  assign {FA_cout_1276,FA_out_1276}=inp_59[54]+inp_60[53]+inp_61[52];
  assign {FA_cout_1277,FA_out_1277}=inp_59[57]+inp_60[56]+inp_61[55];
  assign {FA_cout_1278,FA_out_1278}=inp_59[60]+inp_60[59]+inp_61[58];
  assign {FA_cout_1279,FA_out_1279}=inp_59[63]+inp_60[62]+inp_61[61];
  assign {FA_cout_1280,FA_out_1280}=inp_60[2]+inp_61[1]+inp_62[0];
  assign {FA_cout_1281,FA_out_1281}=inp_60[3]+inp_61[2]+inp_62[1];
  assign {FA_cout_1282,FA_out_1282}=inp_60[4]+inp_61[3]+inp_62[2];
  assign {FA_cout_1283,FA_out_1283}=inp_60[6]+inp_61[5]+inp_62[4];
  assign {FA_cout_1284,FA_out_1284}=inp_60[9]+inp_61[8]+inp_62[7];
  assign {FA_cout_1285,FA_out_1285}=inp_60[12]+inp_61[11]+inp_62[10];
  assign {FA_cout_1286,FA_out_1286}=inp_60[15]+inp_61[14]+inp_62[13];
  assign {FA_cout_1287,FA_out_1287}=inp_60[18]+inp_61[17]+inp_62[16];
  assign {FA_cout_1288,FA_out_1288}=inp_60[21]+inp_61[20]+inp_62[19];
  assign {FA_cout_1289,FA_out_1289}=inp_60[24]+inp_61[23]+inp_62[22];
  assign {FA_cout_1290,FA_out_1290}=inp_60[27]+inp_61[26]+inp_62[25];
  assign {FA_cout_1291,FA_out_1291}=inp_60[30]+inp_61[29]+inp_62[28];
  assign {FA_cout_1292,FA_out_1292}=inp_60[33]+inp_61[32]+inp_62[31];
  assign {FA_cout_1293,FA_out_1293}=inp_60[36]+inp_61[35]+inp_62[34];
  assign {FA_cout_1294,FA_out_1294}=inp_60[39]+inp_61[38]+inp_62[37];
  assign {FA_cout_1295,FA_out_1295}=inp_60[42]+inp_61[41]+inp_62[40];
  assign {FA_cout_1296,FA_out_1296}=inp_60[45]+inp_61[44]+inp_62[43];
  assign {FA_cout_1297,FA_out_1297}=inp_60[48]+inp_61[47]+inp_62[46];
  assign {FA_cout_1298,FA_out_1298}=inp_60[51]+inp_61[50]+inp_62[49];
  assign {FA_cout_1299,FA_out_1299}=inp_60[54]+inp_61[53]+inp_62[52];
  assign {FA_cout_1300,FA_out_1300}=inp_60[57]+inp_61[56]+inp_62[55];
  assign {FA_cout_1301,FA_out_1301}=inp_60[60]+inp_61[59]+inp_62[58];
  assign {FA_cout_1302,FA_out_1302}=inp_60[63]+inp_61[62]+inp_62[61];
  assign {FA_cout_1303,FA_out_1303}=inp_61[6]+inp_62[5]+inp_63[4];
  assign {FA_cout_1304,FA_out_1304}=inp_61[9]+inp_62[8]+inp_63[7];
  assign {FA_cout_1305,FA_out_1305}=inp_61[12]+inp_62[11]+inp_63[10];
  assign {FA_cout_1306,FA_out_1306}=inp_61[15]+inp_62[14]+inp_63[13];
  assign {FA_cout_1307,FA_out_1307}=inp_61[18]+inp_62[17]+inp_63[16];
  assign {FA_cout_1308,FA_out_1308}=inp_61[21]+inp_62[20]+inp_63[19];
  assign {FA_cout_1309,FA_out_1309}=inp_61[24]+inp_62[23]+inp_63[22];
  assign {FA_cout_1310,FA_out_1310}=inp_61[27]+inp_62[26]+inp_63[25];
  assign {FA_cout_1311,FA_out_1311}=inp_61[30]+inp_62[29]+inp_63[28];
  assign {FA_cout_1312,FA_out_1312}=inp_61[33]+inp_62[32]+inp_63[31];
  assign {FA_cout_1313,FA_out_1313}=inp_61[36]+inp_62[35]+inp_63[34];
  assign {FA_cout_1314,FA_out_1314}=inp_61[39]+inp_62[38]+inp_63[37];
  assign {FA_cout_1315,FA_out_1315}=inp_61[42]+inp_62[41]+inp_63[40];
  assign {FA_cout_1316,FA_out_1316}=inp_61[45]+inp_62[44]+inp_63[43];
  assign {FA_cout_1317,FA_out_1317}=inp_61[48]+inp_62[47]+inp_63[46];
  assign {FA_cout_1318,FA_out_1318}=inp_61[51]+inp_62[50]+inp_63[49];
  assign {FA_cout_1319,FA_out_1319}=inp_61[54]+inp_62[53]+inp_63[52];
  assign {FA_cout_1320,FA_out_1320}=inp_61[57]+inp_62[56]+inp_63[55];
  assign {FA_cout_1321,FA_out_1321}=inp_61[60]+inp_62[59]+inp_63[58];
  assign {FA_cout_1322,FA_out_1322}=inp_61[63]+inp_62[62]+inp_63[61];
  assign {FA_cout_1323,FA_out_1323}=FA_cout_0+FA_out_1+inp_3[0];
  assign {FA_cout_1324,FA_out_1324}=FA_cout_1+FA_out_2+HA_out_1;
  assign {FA_cout_1325,FA_out_1325}=FA_cout_2+FA_out_3+HA_cout_1;
  assign {FA_cout_1326,FA_out_1326}=FA_cout_3+FA_out_4+FA_cout_64;
  assign {FA_cout_1327,FA_out_1327}=FA_cout_4+FA_out_5+FA_cout_65;
  assign {FA_cout_1328,FA_out_1328}=FA_cout_5+FA_out_6+FA_cout_66;
  assign {FA_cout_1329,FA_out_1329}=FA_cout_6+FA_out_7+FA_cout_67;
  assign {FA_cout_1330,FA_out_1330}=FA_cout_7+FA_out_8+FA_cout_68;
  assign {FA_cout_1331,FA_out_1331}=FA_cout_8+FA_out_9+FA_cout_69;
  assign {FA_cout_1332,FA_out_1332}=FA_cout_9+FA_out_10+FA_cout_70;
  assign {FA_cout_1333,FA_out_1333}=FA_cout_10+FA_out_11+FA_cout_71;
  assign {FA_cout_1334,FA_out_1334}=FA_cout_11+FA_out_12+FA_cout_72;
  assign {FA_cout_1335,FA_out_1335}=FA_cout_12+FA_out_13+FA_cout_73;
  assign {FA_cout_1336,FA_out_1336}=FA_cout_13+FA_out_14+FA_cout_74;
  assign {FA_cout_1337,FA_out_1337}=FA_cout_14+FA_out_15+FA_cout_75;
  assign {FA_cout_1338,FA_out_1338}=FA_cout_15+FA_out_16+FA_cout_76;
  assign {FA_cout_1339,FA_out_1339}=FA_cout_16+FA_out_17+FA_cout_77;
  assign {FA_cout_1340,FA_out_1340}=FA_cout_17+FA_out_18+FA_cout_78;
  assign {FA_cout_1341,FA_out_1341}=FA_cout_18+FA_out_19+FA_cout_79;
  assign {FA_cout_1342,FA_out_1342}=FA_cout_19+FA_out_20+FA_cout_80;
  assign {FA_cout_1343,FA_out_1343}=FA_cout_20+FA_out_21+FA_cout_81;
  assign {FA_cout_1344,FA_out_1344}=FA_cout_21+FA_out_22+FA_cout_82;
  assign {FA_cout_1345,FA_out_1345}=FA_cout_22+FA_out_23+FA_cout_83;
  assign {FA_cout_1346,FA_out_1346}=FA_cout_23+FA_out_24+FA_cout_84;
  assign {FA_cout_1347,FA_out_1347}=FA_cout_24+FA_out_25+FA_cout_85;
  assign {FA_cout_1348,FA_out_1348}=FA_cout_25+FA_out_26+FA_cout_86;
  assign {FA_cout_1349,FA_out_1349}=FA_cout_26+FA_out_27+FA_cout_87;
  assign {FA_cout_1350,FA_out_1350}=FA_cout_27+FA_out_28+FA_cout_88;
  assign {FA_cout_1351,FA_out_1351}=FA_cout_28+FA_out_29+FA_cout_89;
  assign {FA_cout_1352,FA_out_1352}=FA_cout_29+FA_out_30+FA_cout_90;
  assign {FA_cout_1353,FA_out_1353}=FA_cout_30+FA_out_31+FA_cout_91;
  assign {FA_cout_1354,FA_out_1354}=FA_cout_31+FA_out_32+FA_cout_92;
  assign {FA_cout_1355,FA_out_1355}=FA_cout_32+FA_out_33+FA_cout_93;
  assign {FA_cout_1356,FA_out_1356}=FA_cout_33+FA_out_34+FA_cout_94;
  assign {FA_cout_1357,FA_out_1357}=FA_cout_34+FA_out_35+FA_cout_95;
  assign {FA_cout_1358,FA_out_1358}=FA_cout_35+FA_out_36+FA_cout_96;
  assign {FA_cout_1359,FA_out_1359}=FA_cout_36+FA_out_37+FA_cout_97;
  assign {FA_cout_1360,FA_out_1360}=FA_cout_37+FA_out_38+FA_cout_98;
  assign {FA_cout_1361,FA_out_1361}=FA_cout_38+FA_out_39+FA_cout_99;
  assign {FA_cout_1362,FA_out_1362}=FA_cout_39+FA_out_40+FA_cout_100;
  assign {FA_cout_1363,FA_out_1363}=FA_cout_40+FA_out_41+FA_cout_101;
  assign {FA_cout_1364,FA_out_1364}=FA_cout_41+FA_out_42+FA_cout_102;
  assign {FA_cout_1365,FA_out_1365}=FA_cout_42+FA_out_43+FA_cout_103;
  assign {FA_cout_1366,FA_out_1366}=FA_cout_43+FA_out_44+FA_cout_104;
  assign {FA_cout_1367,FA_out_1367}=FA_cout_44+FA_out_45+FA_cout_105;
  assign {FA_cout_1368,FA_out_1368}=FA_cout_45+FA_out_46+FA_cout_106;
  assign {FA_cout_1369,FA_out_1369}=FA_cout_46+FA_out_47+FA_cout_107;
  assign {FA_cout_1370,FA_out_1370}=FA_cout_47+FA_out_48+FA_cout_108;
  assign {FA_cout_1371,FA_out_1371}=FA_cout_48+FA_out_49+FA_cout_109;
  assign {FA_cout_1372,FA_out_1372}=FA_cout_49+FA_out_50+FA_cout_110;
  assign {FA_cout_1373,FA_out_1373}=FA_cout_50+FA_out_51+FA_cout_111;
  assign {FA_cout_1374,FA_out_1374}=FA_cout_51+FA_out_52+FA_cout_112;
  assign {FA_cout_1375,FA_out_1375}=FA_cout_52+FA_out_53+FA_cout_113;
  assign {FA_cout_1376,FA_out_1376}=FA_cout_53+FA_out_54+FA_cout_114;
  assign {FA_cout_1377,FA_out_1377}=FA_cout_54+FA_out_55+FA_cout_115;
  assign {FA_cout_1378,FA_out_1378}=FA_cout_55+FA_out_56+FA_cout_116;
  assign {FA_cout_1379,FA_out_1379}=FA_cout_56+FA_out_57+FA_cout_117;
  assign {FA_cout_1380,FA_out_1380}=FA_cout_57+FA_out_58+FA_cout_118;
  assign {FA_cout_1381,FA_out_1381}=FA_cout_58+FA_out_59+FA_cout_119;
  assign {FA_cout_1382,FA_out_1382}=FA_cout_59+FA_out_60+FA_cout_120;
  assign {FA_cout_1383,FA_out_1383}=FA_cout_60+FA_out_61+FA_cout_121;
  assign {FA_cout_1384,FA_out_1384}=FA_cout_61+FA_out_62+FA_cout_122;
  assign {FA_cout_1385,FA_out_1385}=FA_cout_62+FA_out_63+FA_cout_123;
  assign {FA_cout_1386,FA_out_1386}=FA_cout_63+FA_out_124+FA_cout_126;
  assign {FA_cout_1387,FA_out_1387}=FA_cout_124+FA_out_125+FA_cout_185;
  assign {FA_cout_1388,FA_out_1388}=FA_out_67+HA_cout_2+FA_out_128;
  assign {FA_cout_1389,FA_out_1389}=FA_out_68+FA_cout_128+FA_out_129;
  assign {FA_cout_1390,FA_out_1390}=FA_out_69+FA_cout_129+FA_out_130;
  assign {FA_cout_1391,FA_out_1391}=FA_out_70+FA_cout_130+FA_out_131;
  assign {FA_cout_1392,FA_out_1392}=FA_out_71+FA_cout_131+FA_out_132;
  assign {FA_cout_1393,FA_out_1393}=FA_out_72+FA_cout_132+FA_out_133;
  assign {FA_cout_1394,FA_out_1394}=FA_out_73+FA_cout_133+FA_out_134;
  assign {FA_cout_1395,FA_out_1395}=FA_out_74+FA_cout_134+FA_out_135;
  assign {FA_cout_1396,FA_out_1396}=FA_out_75+FA_cout_135+FA_out_136;
  assign {FA_cout_1397,FA_out_1397}=FA_out_76+FA_cout_136+FA_out_137;
  assign {FA_cout_1398,FA_out_1398}=FA_out_77+FA_cout_137+FA_out_138;
  assign {FA_cout_1399,FA_out_1399}=FA_out_78+FA_cout_138+FA_out_139;
  assign {FA_cout_1400,FA_out_1400}=FA_out_79+FA_cout_139+FA_out_140;
  assign {FA_cout_1401,FA_out_1401}=FA_out_80+FA_cout_140+FA_out_141;
  assign {FA_cout_1402,FA_out_1402}=FA_out_81+FA_cout_141+FA_out_142;
  assign {FA_cout_1403,FA_out_1403}=FA_out_82+FA_cout_142+FA_out_143;
  assign {FA_cout_1404,FA_out_1404}=FA_out_83+FA_cout_143+FA_out_144;
  assign {FA_cout_1405,FA_out_1405}=FA_out_84+FA_cout_144+FA_out_145;
  assign {FA_cout_1406,FA_out_1406}=FA_out_85+FA_cout_145+FA_out_146;
  assign {FA_cout_1407,FA_out_1407}=FA_out_86+FA_cout_146+FA_out_147;
  assign {FA_cout_1408,FA_out_1408}=FA_out_87+FA_cout_147+FA_out_148;
  assign {FA_cout_1409,FA_out_1409}=FA_out_88+FA_cout_148+FA_out_149;
  assign {FA_cout_1410,FA_out_1410}=FA_out_89+FA_cout_149+FA_out_150;
  assign {FA_cout_1411,FA_out_1411}=FA_out_90+FA_cout_150+FA_out_151;
  assign {FA_cout_1412,FA_out_1412}=FA_out_91+FA_cout_151+FA_out_152;
  assign {FA_cout_1413,FA_out_1413}=FA_out_92+FA_cout_152+FA_out_153;
  assign {FA_cout_1414,FA_out_1414}=FA_out_93+FA_cout_153+FA_out_154;
  assign {FA_cout_1415,FA_out_1415}=FA_out_94+FA_cout_154+FA_out_155;
  assign {FA_cout_1416,FA_out_1416}=FA_out_95+FA_cout_155+FA_out_156;
  assign {FA_cout_1417,FA_out_1417}=FA_out_96+FA_cout_156+FA_out_157;
  assign {FA_cout_1418,FA_out_1418}=FA_out_97+FA_cout_157+FA_out_158;
  assign {FA_cout_1419,FA_out_1419}=FA_out_98+FA_cout_158+FA_out_159;
  assign {FA_cout_1420,FA_out_1420}=FA_out_99+FA_cout_159+FA_out_160;
  assign {FA_cout_1421,FA_out_1421}=FA_out_100+FA_cout_160+FA_out_161;
  assign {FA_cout_1422,FA_out_1422}=FA_out_101+FA_cout_161+FA_out_162;
  assign {FA_cout_1423,FA_out_1423}=FA_out_102+FA_cout_162+FA_out_163;
  assign {FA_cout_1424,FA_out_1424}=FA_out_103+FA_cout_163+FA_out_164;
  assign {FA_cout_1425,FA_out_1425}=FA_out_104+FA_cout_164+FA_out_165;
  assign {FA_cout_1426,FA_out_1426}=FA_out_105+FA_cout_165+FA_out_166;
  assign {FA_cout_1427,FA_out_1427}=FA_out_106+FA_cout_166+FA_out_167;
  assign {FA_cout_1428,FA_out_1428}=FA_out_107+FA_cout_167+FA_out_168;
  assign {FA_cout_1429,FA_out_1429}=FA_out_108+FA_cout_168+FA_out_169;
  assign {FA_cout_1430,FA_out_1430}=FA_out_109+FA_cout_169+FA_out_170;
  assign {FA_cout_1431,FA_out_1431}=FA_out_110+FA_cout_170+FA_out_171;
  assign {FA_cout_1432,FA_out_1432}=FA_out_111+FA_cout_171+FA_out_172;
  assign {FA_cout_1433,FA_out_1433}=FA_out_112+FA_cout_172+FA_out_173;
  assign {FA_cout_1434,FA_out_1434}=FA_out_113+FA_cout_173+FA_out_174;
  assign {FA_cout_1435,FA_out_1435}=FA_out_114+FA_cout_174+FA_out_175;
  assign {FA_cout_1436,FA_out_1436}=FA_out_115+FA_cout_175+FA_out_176;
  assign {FA_cout_1437,FA_out_1437}=FA_out_116+FA_cout_176+FA_out_177;
  assign {FA_cout_1438,FA_out_1438}=FA_out_117+FA_cout_177+FA_out_178;
  assign {FA_cout_1439,FA_out_1439}=FA_out_118+FA_cout_178+FA_out_179;
  assign {FA_cout_1440,FA_out_1440}=FA_out_119+FA_cout_179+FA_out_180;
  assign {FA_cout_1441,FA_out_1441}=FA_out_120+FA_cout_180+FA_out_181;
  assign {FA_cout_1442,FA_out_1442}=FA_out_121+FA_cout_181+FA_out_182;
  assign {FA_cout_1443,FA_out_1443}=FA_out_122+FA_cout_182+FA_out_183;
  assign {FA_cout_1444,FA_out_1444}=FA_out_123+FA_cout_183+FA_out_184;
  assign {FA_cout_1445,FA_out_1445}=FA_cout_125+FA_out_127+FA_cout_187;
  assign {FA_cout_1446,FA_out_1446}=FA_out_126+FA_cout_184+FA_out_189;
  assign {FA_cout_1447,FA_out_1447}=FA_cout_127+FA_out_186+FA_cout_190;
  assign {FA_cout_1448,FA_out_1448}=FA_out_185+FA_cout_189+FA_out_246;
  assign {FA_cout_1449,FA_out_1449}=FA_cout_186+FA_out_188+FA_cout_247;
  assign {FA_cout_1450,FA_out_1450}=FA_out_187+FA_cout_246+FA_out_249;
  assign {FA_cout_1451,FA_out_1451}=FA_cout_188+FA_out_191+FA_cout_250;
  assign {FA_cout_1452,FA_out_1452}=FA_out_190+FA_cout_249+FA_out_253;
  assign {FA_cout_1453,FA_out_1453}=FA_cout_191+FA_out_248+FA_cout_254;
  assign {FA_cout_1454,FA_out_1454}=FA_cout_192+FA_out_193+inp_12[0];
  assign {FA_cout_1455,FA_out_1455}=FA_cout_193+FA_out_194+HA_out_4;
  assign {FA_cout_1456,FA_out_1456}=FA_cout_194+FA_out_195+HA_cout_4;
  assign {FA_cout_1457,FA_out_1457}=FA_cout_195+FA_out_196+FA_cout_256;
  assign {FA_cout_1458,FA_out_1458}=FA_cout_196+FA_out_197+FA_cout_257;
  assign {FA_cout_1459,FA_out_1459}=FA_cout_197+FA_out_198+FA_cout_258;
  assign {FA_cout_1460,FA_out_1460}=FA_cout_198+FA_out_199+FA_cout_259;
  assign {FA_cout_1461,FA_out_1461}=FA_cout_199+FA_out_200+FA_cout_260;
  assign {FA_cout_1462,FA_out_1462}=FA_cout_200+FA_out_201+FA_cout_261;
  assign {FA_cout_1463,FA_out_1463}=FA_cout_201+FA_out_202+FA_cout_262;
  assign {FA_cout_1464,FA_out_1464}=FA_cout_202+FA_out_203+FA_cout_263;
  assign {FA_cout_1465,FA_out_1465}=FA_cout_203+FA_out_204+FA_cout_264;
  assign {FA_cout_1466,FA_out_1466}=FA_cout_204+FA_out_205+FA_cout_265;
  assign {FA_cout_1467,FA_out_1467}=FA_cout_205+FA_out_206+FA_cout_266;
  assign {FA_cout_1468,FA_out_1468}=FA_cout_206+FA_out_207+FA_cout_267;
  assign {FA_cout_1469,FA_out_1469}=FA_cout_207+FA_out_208+FA_cout_268;
  assign {FA_cout_1470,FA_out_1470}=FA_cout_208+FA_out_209+FA_cout_269;
  assign {FA_cout_1471,FA_out_1471}=FA_cout_209+FA_out_210+FA_cout_270;
  assign {FA_cout_1472,FA_out_1472}=FA_cout_210+FA_out_211+FA_cout_271;
  assign {FA_cout_1473,FA_out_1473}=FA_cout_211+FA_out_212+FA_cout_272;
  assign {FA_cout_1474,FA_out_1474}=FA_cout_212+FA_out_213+FA_cout_273;
  assign {FA_cout_1475,FA_out_1475}=FA_cout_213+FA_out_214+FA_cout_274;
  assign {FA_cout_1476,FA_out_1476}=FA_cout_214+FA_out_215+FA_cout_275;
  assign {FA_cout_1477,FA_out_1477}=FA_cout_215+FA_out_216+FA_cout_276;
  assign {FA_cout_1478,FA_out_1478}=FA_cout_216+FA_out_217+FA_cout_277;
  assign {FA_cout_1479,FA_out_1479}=FA_cout_217+FA_out_218+FA_cout_278;
  assign {FA_cout_1480,FA_out_1480}=FA_cout_218+FA_out_219+FA_cout_279;
  assign {FA_cout_1481,FA_out_1481}=FA_cout_219+FA_out_220+FA_cout_280;
  assign {FA_cout_1482,FA_out_1482}=FA_cout_220+FA_out_221+FA_cout_281;
  assign {FA_cout_1483,FA_out_1483}=FA_cout_221+FA_out_222+FA_cout_282;
  assign {FA_cout_1484,FA_out_1484}=FA_cout_222+FA_out_223+FA_cout_283;
  assign {FA_cout_1485,FA_out_1485}=FA_cout_223+FA_out_224+FA_cout_284;
  assign {FA_cout_1486,FA_out_1486}=FA_cout_224+FA_out_225+FA_cout_285;
  assign {FA_cout_1487,FA_out_1487}=FA_cout_225+FA_out_226+FA_cout_286;
  assign {FA_cout_1488,FA_out_1488}=FA_cout_226+FA_out_227+FA_cout_287;
  assign {FA_cout_1489,FA_out_1489}=FA_cout_227+FA_out_228+FA_cout_288;
  assign {FA_cout_1490,FA_out_1490}=FA_cout_228+FA_out_229+FA_cout_289;
  assign {FA_cout_1491,FA_out_1491}=FA_cout_229+FA_out_230+FA_cout_290;
  assign {FA_cout_1492,FA_out_1492}=FA_cout_230+FA_out_231+FA_cout_291;
  assign {FA_cout_1493,FA_out_1493}=FA_cout_231+FA_out_232+FA_cout_292;
  assign {FA_cout_1494,FA_out_1494}=FA_cout_232+FA_out_233+FA_cout_293;
  assign {FA_cout_1495,FA_out_1495}=FA_cout_233+FA_out_234+FA_cout_294;
  assign {FA_cout_1496,FA_out_1496}=FA_cout_234+FA_out_235+FA_cout_295;
  assign {FA_cout_1497,FA_out_1497}=FA_cout_235+FA_out_236+FA_cout_296;
  assign {FA_cout_1498,FA_out_1498}=FA_cout_236+FA_out_237+FA_cout_297;
  assign {FA_cout_1499,FA_out_1499}=FA_cout_237+FA_out_238+FA_cout_298;
  assign {FA_cout_1500,FA_out_1500}=FA_cout_238+FA_out_239+FA_cout_299;
  assign {FA_cout_1501,FA_out_1501}=FA_cout_239+FA_out_240+FA_cout_300;
  assign {FA_cout_1502,FA_out_1502}=FA_cout_240+FA_out_241+FA_cout_301;
  assign {FA_cout_1503,FA_out_1503}=FA_cout_241+FA_out_242+FA_cout_302;
  assign {FA_cout_1504,FA_out_1504}=FA_cout_242+FA_out_243+FA_cout_303;
  assign {FA_cout_1505,FA_out_1505}=FA_cout_243+FA_out_244+FA_cout_304;
  assign {FA_cout_1506,FA_out_1506}=FA_cout_244+FA_out_245+FA_cout_305;
  assign {FA_cout_1507,FA_out_1507}=FA_cout_245+FA_out_252+FA_cout_306;
  assign {FA_cout_1508,FA_out_1508}=FA_out_247+FA_cout_253+FA_out_308;
  assign {FA_cout_1509,FA_out_1509}=FA_cout_248+FA_out_251+FA_cout_309;
  assign {FA_cout_1510,FA_out_1510}=FA_out_250+FA_cout_308+FA_out_312;
  assign {FA_cout_1511,FA_out_1511}=FA_cout_251+FA_out_255+FA_cout_313;
  assign {FA_cout_1512,FA_out_1512}=FA_cout_252+FA_out_307+FA_cout_315;
  assign {FA_cout_1513,FA_out_1513}=FA_out_254+FA_cout_312+FA_out_317;
  assign {FA_cout_1514,FA_out_1514}=FA_cout_255+FA_out_310+FA_cout_318;
  assign {FA_cout_1515,FA_out_1515}=FA_cout_307+FA_out_311+FA_cout_368;
  assign {FA_cout_1516,FA_out_1516}=FA_out_309+FA_cout_317+FA_out_370;
  assign {FA_cout_1517,FA_out_1517}=FA_cout_310+FA_out_314+FA_cout_371;
  assign {FA_cout_1518,FA_out_1518}=FA_out_259+HA_cout_5+FA_out_320;
  assign {FA_cout_1519,FA_out_1519}=FA_out_260+FA_cout_320+FA_out_321;
  assign {FA_cout_1520,FA_out_1520}=FA_out_261+FA_cout_321+FA_out_322;
  assign {FA_cout_1521,FA_out_1521}=FA_out_262+FA_cout_322+FA_out_323;
  assign {FA_cout_1522,FA_out_1522}=FA_out_263+FA_cout_323+FA_out_324;
  assign {FA_cout_1523,FA_out_1523}=FA_out_264+FA_cout_324+FA_out_325;
  assign {FA_cout_1524,FA_out_1524}=FA_out_265+FA_cout_325+FA_out_326;
  assign {FA_cout_1525,FA_out_1525}=FA_out_266+FA_cout_326+FA_out_327;
  assign {FA_cout_1526,FA_out_1526}=FA_out_267+FA_cout_327+FA_out_328;
  assign {FA_cout_1527,FA_out_1527}=FA_out_268+FA_cout_328+FA_out_329;
  assign {FA_cout_1528,FA_out_1528}=FA_out_269+FA_cout_329+FA_out_330;
  assign {FA_cout_1529,FA_out_1529}=FA_out_270+FA_cout_330+FA_out_331;
  assign {FA_cout_1530,FA_out_1530}=FA_out_271+FA_cout_331+FA_out_332;
  assign {FA_cout_1531,FA_out_1531}=FA_out_272+FA_cout_332+FA_out_333;
  assign {FA_cout_1532,FA_out_1532}=FA_out_273+FA_cout_333+FA_out_334;
  assign {FA_cout_1533,FA_out_1533}=FA_out_274+FA_cout_334+FA_out_335;
  assign {FA_cout_1534,FA_out_1534}=FA_out_275+FA_cout_335+FA_out_336;
  assign {FA_cout_1535,FA_out_1535}=FA_out_276+FA_cout_336+FA_out_337;
  assign {FA_cout_1536,FA_out_1536}=FA_out_277+FA_cout_337+FA_out_338;
  assign {FA_cout_1537,FA_out_1537}=FA_out_278+FA_cout_338+FA_out_339;
  assign {FA_cout_1538,FA_out_1538}=FA_out_279+FA_cout_339+FA_out_340;
  assign {FA_cout_1539,FA_out_1539}=FA_out_280+FA_cout_340+FA_out_341;
  assign {FA_cout_1540,FA_out_1540}=FA_out_281+FA_cout_341+FA_out_342;
  assign {FA_cout_1541,FA_out_1541}=FA_out_282+FA_cout_342+FA_out_343;
  assign {FA_cout_1542,FA_out_1542}=FA_out_283+FA_cout_343+FA_out_344;
  assign {FA_cout_1543,FA_out_1543}=FA_out_284+FA_cout_344+FA_out_345;
  assign {FA_cout_1544,FA_out_1544}=FA_out_285+FA_cout_345+FA_out_346;
  assign {FA_cout_1545,FA_out_1545}=FA_out_286+FA_cout_346+FA_out_347;
  assign {FA_cout_1546,FA_out_1546}=FA_out_287+FA_cout_347+FA_out_348;
  assign {FA_cout_1547,FA_out_1547}=FA_out_288+FA_cout_348+FA_out_349;
  assign {FA_cout_1548,FA_out_1548}=FA_out_289+FA_cout_349+FA_out_350;
  assign {FA_cout_1549,FA_out_1549}=FA_out_290+FA_cout_350+FA_out_351;
  assign {FA_cout_1550,FA_out_1550}=FA_out_291+FA_cout_351+FA_out_352;
  assign {FA_cout_1551,FA_out_1551}=FA_out_292+FA_cout_352+FA_out_353;
  assign {FA_cout_1552,FA_out_1552}=FA_out_293+FA_cout_353+FA_out_354;
  assign {FA_cout_1553,FA_out_1553}=FA_out_294+FA_cout_354+FA_out_355;
  assign {FA_cout_1554,FA_out_1554}=FA_out_295+FA_cout_355+FA_out_356;
  assign {FA_cout_1555,FA_out_1555}=FA_out_296+FA_cout_356+FA_out_357;
  assign {FA_cout_1556,FA_out_1556}=FA_out_297+FA_cout_357+FA_out_358;
  assign {FA_cout_1557,FA_out_1557}=FA_out_298+FA_cout_358+FA_out_359;
  assign {FA_cout_1558,FA_out_1558}=FA_out_299+FA_cout_359+FA_out_360;
  assign {FA_cout_1559,FA_out_1559}=FA_out_300+FA_cout_360+FA_out_361;
  assign {FA_cout_1560,FA_out_1560}=FA_out_301+FA_cout_361+FA_out_362;
  assign {FA_cout_1561,FA_out_1561}=FA_out_302+FA_cout_362+FA_out_363;
  assign {FA_cout_1562,FA_out_1562}=FA_out_303+FA_cout_363+FA_out_364;
  assign {FA_cout_1563,FA_out_1563}=FA_out_304+FA_cout_364+FA_out_365;
  assign {FA_cout_1564,FA_out_1564}=FA_out_305+FA_cout_365+FA_out_366;
  assign {FA_cout_1565,FA_out_1565}=FA_out_306+FA_cout_366+FA_out_367;
  assign {FA_cout_1566,FA_out_1566}=FA_cout_311+FA_out_316+FA_cout_373;
  assign {FA_cout_1567,FA_out_1567}=FA_out_313+FA_cout_370+FA_out_375;
  assign {FA_cout_1568,FA_out_1568}=FA_cout_314+FA_out_319+FA_cout_376;
  assign {FA_cout_1569,FA_out_1569}=FA_out_315+FA_cout_367+FA_out_378;
  assign {FA_cout_1570,FA_out_1570}=FA_cout_316+FA_out_369+FA_cout_379;
  assign {FA_cout_1571,FA_out_1571}=FA_out_318+FA_cout_375+FA_out_381;
  assign {FA_cout_1572,FA_out_1572}=FA_cout_319+FA_out_372+FA_cout_382;
  assign {FA_cout_1573,FA_out_1573}=FA_out_368+FA_cout_378+FA_out_429;
  assign {FA_cout_1574,FA_out_1574}=FA_cout_369+FA_out_374+FA_cout_430;
  assign {FA_cout_1575,FA_out_1575}=FA_out_371+FA_cout_381+FA_out_432;
  assign {FA_cout_1576,FA_out_1576}=FA_cout_372+FA_out_377+FA_cout_433;
  assign {FA_cout_1577,FA_out_1577}=FA_out_373+FA_cout_429+FA_out_435;
  assign {FA_cout_1578,FA_out_1578}=FA_cout_374+FA_out_380+FA_cout_436;
  assign {FA_cout_1579,FA_out_1579}=FA_out_376+FA_cout_432+FA_out_438;
  assign {FA_cout_1580,FA_out_1580}=FA_cout_377+FA_out_383+FA_cout_439;
  assign {FA_cout_1581,FA_out_1581}=FA_out_379+FA_cout_435+FA_out_442;
  assign {FA_cout_1582,FA_out_1582}=FA_cout_380+FA_out_431+FA_cout_443;
  assign {FA_cout_1583,FA_out_1583}=FA_out_382+FA_cout_438+FA_out_445;
  assign {FA_cout_1584,FA_out_1584}=FA_cout_383+FA_out_434+FA_cout_446;
  assign {FA_cout_1585,FA_out_1585}=FA_cout_384+FA_out_385+inp_21[0];
  assign {FA_cout_1586,FA_out_1586}=FA_cout_385+FA_out_386+HA_out_7;
  assign {FA_cout_1587,FA_out_1587}=FA_cout_386+FA_out_387+HA_cout_7;
  assign {FA_cout_1588,FA_out_1588}=FA_cout_387+FA_out_388+FA_cout_448;
  assign {FA_cout_1589,FA_out_1589}=FA_cout_388+FA_out_389+FA_cout_449;
  assign {FA_cout_1590,FA_out_1590}=FA_cout_389+FA_out_390+FA_cout_450;
  assign {FA_cout_1591,FA_out_1591}=FA_cout_390+FA_out_391+FA_cout_451;
  assign {FA_cout_1592,FA_out_1592}=FA_cout_391+FA_out_392+FA_cout_452;
  assign {FA_cout_1593,FA_out_1593}=FA_cout_392+FA_out_393+FA_cout_453;
  assign {FA_cout_1594,FA_out_1594}=FA_cout_393+FA_out_394+FA_cout_454;
  assign {FA_cout_1595,FA_out_1595}=FA_cout_394+FA_out_395+FA_cout_455;
  assign {FA_cout_1596,FA_out_1596}=FA_cout_395+FA_out_396+FA_cout_456;
  assign {FA_cout_1597,FA_out_1597}=FA_cout_396+FA_out_397+FA_cout_457;
  assign {FA_cout_1598,FA_out_1598}=FA_cout_397+FA_out_398+FA_cout_458;
  assign {FA_cout_1599,FA_out_1599}=FA_cout_398+FA_out_399+FA_cout_459;
  assign {FA_cout_1600,FA_out_1600}=FA_cout_399+FA_out_400+FA_cout_460;
  assign {FA_cout_1601,FA_out_1601}=FA_cout_400+FA_out_401+FA_cout_461;
  assign {FA_cout_1602,FA_out_1602}=FA_cout_401+FA_out_402+FA_cout_462;
  assign {FA_cout_1603,FA_out_1603}=FA_cout_402+FA_out_403+FA_cout_463;
  assign {FA_cout_1604,FA_out_1604}=FA_cout_403+FA_out_404+FA_cout_464;
  assign {FA_cout_1605,FA_out_1605}=FA_cout_404+FA_out_405+FA_cout_465;
  assign {FA_cout_1606,FA_out_1606}=FA_cout_405+FA_out_406+FA_cout_466;
  assign {FA_cout_1607,FA_out_1607}=FA_cout_406+FA_out_407+FA_cout_467;
  assign {FA_cout_1608,FA_out_1608}=FA_cout_407+FA_out_408+FA_cout_468;
  assign {FA_cout_1609,FA_out_1609}=FA_cout_408+FA_out_409+FA_cout_469;
  assign {FA_cout_1610,FA_out_1610}=FA_cout_409+FA_out_410+FA_cout_470;
  assign {FA_cout_1611,FA_out_1611}=FA_cout_410+FA_out_411+FA_cout_471;
  assign {FA_cout_1612,FA_out_1612}=FA_cout_411+FA_out_412+FA_cout_472;
  assign {FA_cout_1613,FA_out_1613}=FA_cout_412+FA_out_413+FA_cout_473;
  assign {FA_cout_1614,FA_out_1614}=FA_cout_413+FA_out_414+FA_cout_474;
  assign {FA_cout_1615,FA_out_1615}=FA_cout_414+FA_out_415+FA_cout_475;
  assign {FA_cout_1616,FA_out_1616}=FA_cout_415+FA_out_416+FA_cout_476;
  assign {FA_cout_1617,FA_out_1617}=FA_cout_416+FA_out_417+FA_cout_477;
  assign {FA_cout_1618,FA_out_1618}=FA_cout_417+FA_out_418+FA_cout_478;
  assign {FA_cout_1619,FA_out_1619}=FA_cout_418+FA_out_419+FA_cout_479;
  assign {FA_cout_1620,FA_out_1620}=FA_cout_419+FA_out_420+FA_cout_480;
  assign {FA_cout_1621,FA_out_1621}=FA_cout_420+FA_out_421+FA_cout_481;
  assign {FA_cout_1622,FA_out_1622}=FA_cout_421+FA_out_422+FA_cout_482;
  assign {FA_cout_1623,FA_out_1623}=FA_cout_422+FA_out_423+FA_cout_483;
  assign {FA_cout_1624,FA_out_1624}=FA_cout_423+FA_out_424+FA_cout_484;
  assign {FA_cout_1625,FA_out_1625}=FA_cout_424+FA_out_425+FA_cout_485;
  assign {FA_cout_1626,FA_out_1626}=FA_cout_425+FA_out_426+FA_cout_486;
  assign {FA_cout_1627,FA_out_1627}=FA_cout_426+FA_out_427+FA_cout_487;
  assign {FA_cout_1628,FA_out_1628}=FA_cout_427+FA_out_428+FA_cout_488;
  assign {FA_cout_1629,FA_out_1629}=FA_cout_428+FA_out_441+FA_cout_489;
  assign {FA_cout_1630,FA_out_1630}=FA_out_430+FA_cout_442+FA_out_491;
  assign {FA_cout_1631,FA_out_1631}=FA_cout_431+FA_out_437+FA_cout_492;
  assign {FA_cout_1632,FA_out_1632}=FA_out_433+FA_cout_445+FA_out_494;
  assign {FA_cout_1633,FA_out_1633}=FA_cout_434+FA_out_440+FA_cout_495;
  assign {FA_cout_1634,FA_out_1634}=FA_out_436+FA_cout_491+FA_out_498;
  assign {FA_cout_1635,FA_out_1635}=FA_cout_437+FA_out_444+FA_cout_499;
  assign {FA_cout_1636,FA_out_1636}=FA_out_439+FA_cout_494+FA_out_501;
  assign {FA_cout_1637,FA_out_1637}=FA_cout_440+FA_out_447+FA_cout_502;
  assign {FA_cout_1638,FA_out_1638}=FA_cout_441+FA_out_490+FA_cout_504;
  assign {FA_cout_1639,FA_out_1639}=FA_out_443+FA_cout_498+FA_out_506;
  assign {FA_cout_1640,FA_out_1640}=FA_cout_444+FA_out_493+FA_cout_507;
  assign {FA_cout_1641,FA_out_1641}=FA_out_446+FA_cout_501+FA_out_509;
  assign {FA_cout_1642,FA_out_1642}=FA_cout_447+FA_out_496+FA_cout_510;
  assign {FA_cout_1643,FA_out_1643}=FA_cout_490+FA_out_497+FA_cout_551;
  assign {FA_cout_1644,FA_out_1644}=FA_out_492+FA_cout_506+FA_out_553;
  assign {FA_cout_1645,FA_out_1645}=FA_cout_493+FA_out_500+FA_cout_554;
  assign {FA_cout_1646,FA_out_1646}=FA_out_495+FA_cout_509+FA_out_556;
  assign {FA_cout_1647,FA_out_1647}=FA_cout_496+FA_out_503+FA_cout_557;
  assign {FA_cout_1648,FA_out_1648}=FA_out_451+HA_cout_8+FA_out_512;
  assign {FA_cout_1649,FA_out_1649}=FA_out_452+FA_cout_512+FA_out_513;
  assign {FA_cout_1650,FA_out_1650}=FA_out_453+FA_cout_513+FA_out_514;
  assign {FA_cout_1651,FA_out_1651}=FA_out_454+FA_cout_514+FA_out_515;
  assign {FA_cout_1652,FA_out_1652}=FA_out_455+FA_cout_515+FA_out_516;
  assign {FA_cout_1653,FA_out_1653}=FA_out_456+FA_cout_516+FA_out_517;
  assign {FA_cout_1654,FA_out_1654}=FA_out_457+FA_cout_517+FA_out_518;
  assign {FA_cout_1655,FA_out_1655}=FA_out_458+FA_cout_518+FA_out_519;
  assign {FA_cout_1656,FA_out_1656}=FA_out_459+FA_cout_519+FA_out_520;
  assign {FA_cout_1657,FA_out_1657}=FA_out_460+FA_cout_520+FA_out_521;
  assign {FA_cout_1658,FA_out_1658}=FA_out_461+FA_cout_521+FA_out_522;
  assign {FA_cout_1659,FA_out_1659}=FA_out_462+FA_cout_522+FA_out_523;
  assign {FA_cout_1660,FA_out_1660}=FA_out_463+FA_cout_523+FA_out_524;
  assign {FA_cout_1661,FA_out_1661}=FA_out_464+FA_cout_524+FA_out_525;
  assign {FA_cout_1662,FA_out_1662}=FA_out_465+FA_cout_525+FA_out_526;
  assign {FA_cout_1663,FA_out_1663}=FA_out_466+FA_cout_526+FA_out_527;
  assign {FA_cout_1664,FA_out_1664}=FA_out_467+FA_cout_527+FA_out_528;
  assign {FA_cout_1665,FA_out_1665}=FA_out_468+FA_cout_528+FA_out_529;
  assign {FA_cout_1666,FA_out_1666}=FA_out_469+FA_cout_529+FA_out_530;
  assign {FA_cout_1667,FA_out_1667}=FA_out_470+FA_cout_530+FA_out_531;
  assign {FA_cout_1668,FA_out_1668}=FA_out_471+FA_cout_531+FA_out_532;
  assign {FA_cout_1669,FA_out_1669}=FA_out_472+FA_cout_532+FA_out_533;
  assign {FA_cout_1670,FA_out_1670}=FA_out_473+FA_cout_533+FA_out_534;
  assign {FA_cout_1671,FA_out_1671}=FA_out_474+FA_cout_534+FA_out_535;
  assign {FA_cout_1672,FA_out_1672}=FA_out_475+FA_cout_535+FA_out_536;
  assign {FA_cout_1673,FA_out_1673}=FA_out_476+FA_cout_536+FA_out_537;
  assign {FA_cout_1674,FA_out_1674}=FA_out_477+FA_cout_537+FA_out_538;
  assign {FA_cout_1675,FA_out_1675}=FA_out_478+FA_cout_538+FA_out_539;
  assign {FA_cout_1676,FA_out_1676}=FA_out_479+FA_cout_539+FA_out_540;
  assign {FA_cout_1677,FA_out_1677}=FA_out_480+FA_cout_540+FA_out_541;
  assign {FA_cout_1678,FA_out_1678}=FA_out_481+FA_cout_541+FA_out_542;
  assign {FA_cout_1679,FA_out_1679}=FA_out_482+FA_cout_542+FA_out_543;
  assign {FA_cout_1680,FA_out_1680}=FA_out_483+FA_cout_543+FA_out_544;
  assign {FA_cout_1681,FA_out_1681}=FA_out_484+FA_cout_544+FA_out_545;
  assign {FA_cout_1682,FA_out_1682}=FA_out_485+FA_cout_545+FA_out_546;
  assign {FA_cout_1683,FA_out_1683}=FA_out_486+FA_cout_546+FA_out_547;
  assign {FA_cout_1684,FA_out_1684}=FA_out_487+FA_cout_547+FA_out_548;
  assign {FA_cout_1685,FA_out_1685}=FA_out_488+FA_cout_548+FA_out_549;
  assign {FA_cout_1686,FA_out_1686}=FA_out_489+FA_cout_549+FA_out_550;
  assign {FA_cout_1687,FA_out_1687}=FA_cout_497+FA_out_505+FA_cout_559;
  assign {FA_cout_1688,FA_out_1688}=FA_out_499+FA_cout_553+FA_out_561;
  assign {FA_cout_1689,FA_out_1689}=FA_cout_500+FA_out_508+FA_cout_562;
  assign {FA_cout_1690,FA_out_1690}=FA_out_502+FA_cout_556+FA_out_564;
  assign {FA_cout_1691,FA_out_1691}=FA_cout_503+FA_out_511+FA_cout_565;
  assign {FA_cout_1692,FA_out_1692}=FA_out_504+FA_cout_550+FA_out_567;
  assign {FA_cout_1693,FA_out_1693}=FA_cout_505+FA_out_552+FA_cout_568;
  assign {FA_cout_1694,FA_out_1694}=FA_out_507+FA_cout_561+FA_out_570;
  assign {FA_cout_1695,FA_out_1695}=FA_cout_508+FA_out_555+FA_cout_571;
  assign {FA_cout_1696,FA_out_1696}=FA_out_510+FA_cout_564+FA_out_573;
  assign {FA_cout_1697,FA_out_1697}=FA_cout_511+FA_out_558+FA_cout_574;
  assign {FA_cout_1698,FA_out_1698}=FA_out_551+FA_cout_567+FA_out_612;
  assign {FA_cout_1699,FA_out_1699}=FA_cout_552+FA_out_560+FA_cout_613;
  assign {FA_cout_1700,FA_out_1700}=FA_out_554+FA_cout_570+FA_out_615;
  assign {FA_cout_1701,FA_out_1701}=FA_cout_555+FA_out_563+FA_cout_616;
  assign {FA_cout_1702,FA_out_1702}=FA_out_557+FA_cout_573+FA_out_618;
  assign {FA_cout_1703,FA_out_1703}=FA_cout_558+FA_out_566+FA_cout_619;
  assign {FA_cout_1704,FA_out_1704}=FA_out_559+FA_cout_612+FA_out_621;
  assign {FA_cout_1705,FA_out_1705}=FA_cout_560+FA_out_569+FA_cout_622;
  assign {FA_cout_1706,FA_out_1706}=FA_out_562+FA_cout_615+FA_out_624;
  assign {FA_cout_1707,FA_out_1707}=FA_cout_563+FA_out_572+FA_cout_625;
  assign {FA_cout_1708,FA_out_1708}=FA_out_565+FA_cout_618+FA_out_627;
  assign {FA_cout_1709,FA_out_1709}=FA_cout_566+FA_out_575+FA_cout_628;
  assign {FA_cout_1710,FA_out_1710}=FA_out_568+FA_cout_621+FA_out_631;
  assign {FA_cout_1711,FA_out_1711}=FA_cout_569+FA_out_614+FA_cout_632;
  assign {FA_cout_1712,FA_out_1712}=FA_out_571+FA_cout_624+FA_out_634;
  assign {FA_cout_1713,FA_out_1713}=FA_cout_572+FA_out_617+FA_cout_635;
  assign {FA_cout_1714,FA_out_1714}=FA_out_574+FA_cout_627+FA_out_637;
  assign {FA_cout_1715,FA_out_1715}=FA_cout_575+FA_out_620+FA_cout_638;
  assign {FA_cout_1716,FA_out_1716}=FA_cout_576+FA_out_577+inp_30[0];
  assign {FA_cout_1717,FA_out_1717}=FA_cout_577+FA_out_578+HA_out_10;
  assign {FA_cout_1718,FA_out_1718}=FA_cout_578+FA_out_579+HA_cout_10;
  assign {FA_cout_1719,FA_out_1719}=FA_cout_579+FA_out_580+FA_cout_640;
  assign {FA_cout_1720,FA_out_1720}=FA_cout_580+FA_out_581+FA_cout_641;
  assign {FA_cout_1721,FA_out_1721}=FA_cout_581+FA_out_582+FA_cout_642;
  assign {FA_cout_1722,FA_out_1722}=FA_cout_582+FA_out_583+FA_cout_643;
  assign {FA_cout_1723,FA_out_1723}=FA_cout_583+FA_out_584+FA_cout_644;
  assign {FA_cout_1724,FA_out_1724}=FA_cout_584+FA_out_585+FA_cout_645;
  assign {FA_cout_1725,FA_out_1725}=FA_cout_585+FA_out_586+FA_cout_646;
  assign {FA_cout_1726,FA_out_1726}=FA_cout_586+FA_out_587+FA_cout_647;
  assign {FA_cout_1727,FA_out_1727}=FA_cout_587+FA_out_588+FA_cout_648;
  assign {FA_cout_1728,FA_out_1728}=FA_cout_588+FA_out_589+FA_cout_649;
  assign {FA_cout_1729,FA_out_1729}=FA_cout_589+FA_out_590+FA_cout_650;
  assign {FA_cout_1730,FA_out_1730}=FA_cout_590+FA_out_591+FA_cout_651;
  assign {FA_cout_1731,FA_out_1731}=FA_cout_591+FA_out_592+FA_cout_652;
  assign {FA_cout_1732,FA_out_1732}=FA_cout_592+FA_out_593+FA_cout_653;
  assign {FA_cout_1733,FA_out_1733}=FA_cout_593+FA_out_594+FA_cout_654;
  assign {FA_cout_1734,FA_out_1734}=FA_cout_594+FA_out_595+FA_cout_655;
  assign {FA_cout_1735,FA_out_1735}=FA_cout_595+FA_out_596+FA_cout_656;
  assign {FA_cout_1736,FA_out_1736}=FA_cout_596+FA_out_597+FA_cout_657;
  assign {FA_cout_1737,FA_out_1737}=FA_cout_597+FA_out_598+FA_cout_658;
  assign {FA_cout_1738,FA_out_1738}=FA_cout_598+FA_out_599+FA_cout_659;
  assign {FA_cout_1739,FA_out_1739}=FA_cout_599+FA_out_600+FA_cout_660;
  assign {FA_cout_1740,FA_out_1740}=FA_cout_600+FA_out_601+FA_cout_661;
  assign {FA_cout_1741,FA_out_1741}=FA_cout_601+FA_out_602+FA_cout_662;
  assign {FA_cout_1742,FA_out_1742}=FA_cout_602+FA_out_603+FA_cout_663;
  assign {FA_cout_1743,FA_out_1743}=FA_cout_603+FA_out_604+FA_cout_664;
  assign {FA_cout_1744,FA_out_1744}=FA_cout_604+FA_out_605+FA_cout_665;
  assign {FA_cout_1745,FA_out_1745}=FA_cout_605+FA_out_606+FA_cout_666;
  assign {FA_cout_1746,FA_out_1746}=FA_cout_606+FA_out_607+FA_cout_667;
  assign {FA_cout_1747,FA_out_1747}=FA_cout_607+FA_out_608+FA_cout_668;
  assign {FA_cout_1748,FA_out_1748}=FA_cout_608+FA_out_609+FA_cout_669;
  assign {FA_cout_1749,FA_out_1749}=FA_cout_609+FA_out_610+FA_cout_670;
  assign {FA_cout_1750,FA_out_1750}=FA_cout_610+FA_out_611+FA_cout_671;
  assign {FA_cout_1751,FA_out_1751}=FA_cout_611+FA_out_630+FA_cout_672;
  assign {FA_cout_1752,FA_out_1752}=FA_out_613+FA_cout_631+FA_out_674;
  assign {FA_cout_1753,FA_out_1753}=FA_cout_614+FA_out_623+FA_cout_675;
  assign {FA_cout_1754,FA_out_1754}=FA_out_616+FA_cout_634+FA_out_677;
  assign {FA_cout_1755,FA_out_1755}=FA_cout_617+FA_out_626+FA_cout_678;
  assign {FA_cout_1756,FA_out_1756}=FA_out_619+FA_cout_637+FA_out_680;
  assign {FA_cout_1757,FA_out_1757}=FA_cout_620+FA_out_629+FA_cout_681;
  assign {FA_cout_1758,FA_out_1758}=FA_out_622+FA_cout_674+FA_out_684;
  assign {FA_cout_1759,FA_out_1759}=FA_cout_623+FA_out_633+FA_cout_685;
  assign {FA_cout_1760,FA_out_1760}=FA_out_625+FA_cout_677+FA_out_687;
  assign {FA_cout_1761,FA_out_1761}=FA_cout_626+FA_out_636+FA_cout_688;
  assign {FA_cout_1762,FA_out_1762}=FA_out_628+FA_cout_680+FA_out_690;
  assign {FA_cout_1763,FA_out_1763}=FA_cout_629+FA_out_639+FA_cout_691;
  assign {FA_cout_1764,FA_out_1764}=FA_cout_630+FA_out_673+FA_cout_693;
  assign {FA_cout_1765,FA_out_1765}=FA_out_632+FA_cout_684+FA_out_695;
  assign {FA_cout_1766,FA_out_1766}=FA_cout_633+FA_out_676+FA_cout_696;
  assign {FA_cout_1767,FA_out_1767}=FA_out_635+FA_cout_687+FA_out_698;
  assign {FA_cout_1768,FA_out_1768}=FA_cout_636+FA_out_679+FA_cout_699;
  assign {FA_cout_1769,FA_out_1769}=FA_out_638+FA_cout_690+FA_out_701;
  assign {FA_cout_1770,FA_out_1770}=FA_cout_639+FA_out_682+FA_cout_702;
  assign {FA_cout_1771,FA_out_1771}=FA_cout_673+FA_out_683+FA_cout_734;
  assign {FA_cout_1772,FA_out_1772}=FA_out_675+FA_cout_695+FA_out_736;
  assign {FA_cout_1773,FA_out_1773}=FA_cout_676+FA_out_686+FA_cout_737;
  assign {FA_cout_1774,FA_out_1774}=FA_out_678+FA_cout_698+FA_out_739;
  assign {FA_cout_1775,FA_out_1775}=FA_cout_679+FA_out_689+FA_cout_740;
  assign {FA_cout_1776,FA_out_1776}=FA_out_681+FA_cout_701+FA_out_742;
  assign {FA_cout_1777,FA_out_1777}=FA_cout_682+FA_out_692+FA_cout_743;
  assign {FA_cout_1778,FA_out_1778}=FA_out_643+HA_cout_11+FA_out_704;
  assign {FA_cout_1779,FA_out_1779}=FA_out_644+FA_cout_704+FA_out_705;
  assign {FA_cout_1780,FA_out_1780}=FA_out_645+FA_cout_705+FA_out_706;
  assign {FA_cout_1781,FA_out_1781}=FA_out_646+FA_cout_706+FA_out_707;
  assign {FA_cout_1782,FA_out_1782}=FA_out_647+FA_cout_707+FA_out_708;
  assign {FA_cout_1783,FA_out_1783}=FA_out_648+FA_cout_708+FA_out_709;
  assign {FA_cout_1784,FA_out_1784}=FA_out_649+FA_cout_709+FA_out_710;
  assign {FA_cout_1785,FA_out_1785}=FA_out_650+FA_cout_710+FA_out_711;
  assign {FA_cout_1786,FA_out_1786}=FA_out_651+FA_cout_711+FA_out_712;
  assign {FA_cout_1787,FA_out_1787}=FA_out_652+FA_cout_712+FA_out_713;
  assign {FA_cout_1788,FA_out_1788}=FA_out_653+FA_cout_713+FA_out_714;
  assign {FA_cout_1789,FA_out_1789}=FA_out_654+FA_cout_714+FA_out_715;
  assign {FA_cout_1790,FA_out_1790}=FA_out_655+FA_cout_715+FA_out_716;
  assign {FA_cout_1791,FA_out_1791}=FA_out_656+FA_cout_716+FA_out_717;
  assign {FA_cout_1792,FA_out_1792}=FA_out_657+FA_cout_717+FA_out_718;
  assign {FA_cout_1793,FA_out_1793}=FA_out_658+FA_cout_718+FA_out_719;
  assign {FA_cout_1794,FA_out_1794}=FA_out_659+FA_cout_719+FA_out_720;
  assign {FA_cout_1795,FA_out_1795}=FA_out_660+FA_cout_720+FA_out_721;
  assign {FA_cout_1796,FA_out_1796}=FA_out_661+FA_cout_721+FA_out_722;
  assign {FA_cout_1797,FA_out_1797}=FA_out_662+FA_cout_722+FA_out_723;
  assign {FA_cout_1798,FA_out_1798}=FA_out_663+FA_cout_723+FA_out_724;
  assign {FA_cout_1799,FA_out_1799}=FA_out_664+FA_cout_724+FA_out_725;
  assign {FA_cout_1800,FA_out_1800}=FA_out_665+FA_cout_725+FA_out_726;
  assign {FA_cout_1801,FA_out_1801}=FA_out_666+FA_cout_726+FA_out_727;
  assign {FA_cout_1802,FA_out_1802}=FA_out_667+FA_cout_727+FA_out_728;
  assign {FA_cout_1803,FA_out_1803}=FA_out_668+FA_cout_728+FA_out_729;
  assign {FA_cout_1804,FA_out_1804}=FA_out_669+FA_cout_729+FA_out_730;
  assign {FA_cout_1805,FA_out_1805}=FA_out_670+FA_cout_730+FA_out_731;
  assign {FA_cout_1806,FA_out_1806}=FA_out_671+FA_cout_731+FA_out_732;
  assign {FA_cout_1807,FA_out_1807}=FA_out_672+FA_cout_732+FA_out_733;
  assign {FA_cout_1808,FA_out_1808}=FA_cout_683+FA_out_694+FA_cout_745;
  assign {FA_cout_1809,FA_out_1809}=FA_out_685+FA_cout_736+FA_out_747;
  assign {FA_cout_1810,FA_out_1810}=FA_cout_686+FA_out_697+FA_cout_748;
  assign {FA_cout_1811,FA_out_1811}=FA_out_688+FA_cout_739+FA_out_750;
  assign {FA_cout_1812,FA_out_1812}=FA_cout_689+FA_out_700+FA_cout_751;
  assign {FA_cout_1813,FA_out_1813}=FA_out_691+FA_cout_742+FA_out_753;
  assign {FA_cout_1814,FA_out_1814}=FA_cout_692+FA_out_703+FA_cout_754;
  assign {FA_cout_1815,FA_out_1815}=FA_out_693+FA_cout_733+FA_out_756;
  assign {FA_cout_1816,FA_out_1816}=FA_cout_694+FA_out_735+FA_cout_757;
  assign {FA_cout_1817,FA_out_1817}=FA_out_696+FA_cout_747+FA_out_759;
  assign {FA_cout_1818,FA_out_1818}=FA_cout_697+FA_out_738+FA_cout_760;
  assign {FA_cout_1819,FA_out_1819}=FA_out_699+FA_cout_750+FA_out_762;
  assign {FA_cout_1820,FA_out_1820}=FA_cout_700+FA_out_741+FA_cout_763;
  assign {FA_cout_1821,FA_out_1821}=FA_out_702+FA_cout_753+FA_out_765;
  assign {FA_cout_1822,FA_out_1822}=FA_cout_703+FA_out_744+FA_cout_766;
  assign {FA_cout_1823,FA_out_1823}=FA_out_734+FA_cout_756+FA_out_795;
  assign {FA_cout_1824,FA_out_1824}=FA_cout_735+FA_out_746+FA_cout_796;
  assign {FA_cout_1825,FA_out_1825}=FA_out_737+FA_cout_759+FA_out_798;
  assign {FA_cout_1826,FA_out_1826}=FA_cout_738+FA_out_749+FA_cout_799;
  assign {FA_cout_1827,FA_out_1827}=FA_out_740+FA_cout_762+FA_out_801;
  assign {FA_cout_1828,FA_out_1828}=FA_cout_741+FA_out_752+FA_cout_802;
  assign {FA_cout_1829,FA_out_1829}=FA_out_743+FA_cout_765+FA_out_804;
  assign {FA_cout_1830,FA_out_1830}=FA_cout_744+FA_out_755+FA_cout_805;
  assign {FA_cout_1831,FA_out_1831}=FA_out_745+FA_cout_795+FA_out_807;
  assign {FA_cout_1832,FA_out_1832}=FA_cout_746+FA_out_758+FA_cout_808;
  assign {FA_cout_1833,FA_out_1833}=FA_out_748+FA_cout_798+FA_out_810;
  assign {FA_cout_1834,FA_out_1834}=FA_cout_749+FA_out_761+FA_cout_811;
  assign {FA_cout_1835,FA_out_1835}=FA_out_751+FA_cout_801+FA_out_813;
  assign {FA_cout_1836,FA_out_1836}=FA_cout_752+FA_out_764+FA_cout_814;
  assign {FA_cout_1837,FA_out_1837}=FA_out_754+FA_cout_804+FA_out_816;
  assign {FA_cout_1838,FA_out_1838}=FA_cout_755+FA_out_767+FA_cout_817;
  assign {FA_cout_1839,FA_out_1839}=FA_out_757+FA_cout_807+FA_out_820;
  assign {FA_cout_1840,FA_out_1840}=FA_cout_758+FA_out_797+FA_cout_821;
  assign {FA_cout_1841,FA_out_1841}=FA_out_760+FA_cout_810+FA_out_823;
  assign {FA_cout_1842,FA_out_1842}=FA_cout_761+FA_out_800+FA_cout_824;
  assign {FA_cout_1843,FA_out_1843}=FA_out_763+FA_cout_813+FA_out_826;
  assign {FA_cout_1844,FA_out_1844}=FA_cout_764+FA_out_803+FA_cout_827;
  assign {FA_cout_1845,FA_out_1845}=FA_out_766+FA_cout_816+FA_out_829;
  assign {FA_cout_1846,FA_out_1846}=FA_cout_767+FA_out_806+FA_cout_830;
  assign {FA_cout_1847,FA_out_1847}=FA_cout_768+FA_out_769+inp_39[0];
  assign {FA_cout_1848,FA_out_1848}=FA_cout_769+FA_out_770+HA_out_13;
  assign {FA_cout_1849,FA_out_1849}=FA_cout_770+FA_out_771+HA_cout_13;
  assign {FA_cout_1850,FA_out_1850}=FA_cout_771+FA_out_772+FA_cout_832;
  assign {FA_cout_1851,FA_out_1851}=FA_cout_772+FA_out_773+FA_cout_833;
  assign {FA_cout_1852,FA_out_1852}=FA_cout_773+FA_out_774+FA_cout_834;
  assign {FA_cout_1853,FA_out_1853}=FA_cout_774+FA_out_775+FA_cout_835;
  assign {FA_cout_1854,FA_out_1854}=FA_cout_775+FA_out_776+FA_cout_836;
  assign {FA_cout_1855,FA_out_1855}=FA_cout_776+FA_out_777+FA_cout_837;
  assign {FA_cout_1856,FA_out_1856}=FA_cout_777+FA_out_778+FA_cout_838;
  assign {FA_cout_1857,FA_out_1857}=FA_cout_778+FA_out_779+FA_cout_839;
  assign {FA_cout_1858,FA_out_1858}=FA_cout_779+FA_out_780+FA_cout_840;
  assign {FA_cout_1859,FA_out_1859}=FA_cout_780+FA_out_781+FA_cout_841;
  assign {FA_cout_1860,FA_out_1860}=FA_cout_781+FA_out_782+FA_cout_842;
  assign {FA_cout_1861,FA_out_1861}=FA_cout_782+FA_out_783+FA_cout_843;
  assign {FA_cout_1862,FA_out_1862}=FA_cout_783+FA_out_784+FA_cout_844;
  assign {FA_cout_1863,FA_out_1863}=FA_cout_784+FA_out_785+FA_cout_845;
  assign {FA_cout_1864,FA_out_1864}=FA_cout_785+FA_out_786+FA_cout_846;
  assign {FA_cout_1865,FA_out_1865}=FA_cout_786+FA_out_787+FA_cout_847;
  assign {FA_cout_1866,FA_out_1866}=FA_cout_787+FA_out_788+FA_cout_848;
  assign {FA_cout_1867,FA_out_1867}=FA_cout_788+FA_out_789+FA_cout_849;
  assign {FA_cout_1868,FA_out_1868}=FA_cout_789+FA_out_790+FA_cout_850;
  assign {FA_cout_1869,FA_out_1869}=FA_cout_790+FA_out_791+FA_cout_851;
  assign {FA_cout_1870,FA_out_1870}=FA_cout_791+FA_out_792+FA_cout_852;
  assign {FA_cout_1871,FA_out_1871}=FA_cout_792+FA_out_793+FA_cout_853;
  assign {FA_cout_1872,FA_out_1872}=FA_cout_793+FA_out_794+FA_cout_854;
  assign {FA_cout_1873,FA_out_1873}=FA_cout_794+FA_out_819+FA_cout_855;
  assign {FA_cout_1874,FA_out_1874}=FA_out_796+FA_cout_820+FA_out_857;
  assign {FA_cout_1875,FA_out_1875}=FA_cout_797+FA_out_809+FA_cout_858;
  assign {FA_cout_1876,FA_out_1876}=FA_out_799+FA_cout_823+FA_out_860;
  assign {FA_cout_1877,FA_out_1877}=FA_cout_800+FA_out_812+FA_cout_861;
  assign {FA_cout_1878,FA_out_1878}=FA_out_802+FA_cout_826+FA_out_863;
  assign {FA_cout_1879,FA_out_1879}=FA_cout_803+FA_out_815+FA_cout_864;
  assign {FA_cout_1880,FA_out_1880}=FA_out_805+FA_cout_829+FA_out_866;
  assign {FA_cout_1881,FA_out_1881}=FA_cout_806+FA_out_818+FA_cout_867;
  assign {FA_cout_1882,FA_out_1882}=FA_out_808+FA_cout_857+FA_out_870;
  assign {FA_cout_1883,FA_out_1883}=FA_cout_809+FA_out_822+FA_cout_871;
  assign {FA_cout_1884,FA_out_1884}=FA_out_811+FA_cout_860+FA_out_873;
  assign {FA_cout_1885,FA_out_1885}=FA_cout_812+FA_out_825+FA_cout_874;
  assign {FA_cout_1886,FA_out_1886}=FA_out_814+FA_cout_863+FA_out_876;
  assign {FA_cout_1887,FA_out_1887}=FA_cout_815+FA_out_828+FA_cout_877;
  assign {FA_cout_1888,FA_out_1888}=FA_out_817+FA_cout_866+FA_out_879;
  assign {FA_cout_1889,FA_out_1889}=FA_cout_818+FA_out_831+FA_cout_880;
  assign {FA_cout_1890,FA_out_1890}=FA_cout_819+FA_out_856+FA_cout_882;
  assign {FA_cout_1891,FA_out_1891}=FA_out_821+FA_cout_870+FA_out_884;
  assign {FA_cout_1892,FA_out_1892}=FA_cout_822+FA_out_859+FA_cout_885;
  assign {FA_cout_1893,FA_out_1893}=FA_out_824+FA_cout_873+FA_out_887;
  assign {FA_cout_1894,FA_out_1894}=FA_cout_825+FA_out_862+FA_cout_888;
  assign {FA_cout_1895,FA_out_1895}=FA_out_827+FA_cout_876+FA_out_890;
  assign {FA_cout_1896,FA_out_1896}=FA_cout_828+FA_out_865+FA_cout_891;
  assign {FA_cout_1897,FA_out_1897}=FA_out_830+FA_cout_879+FA_out_893;
  assign {FA_cout_1898,FA_out_1898}=FA_cout_831+FA_out_868+FA_cout_894;
  assign {FA_cout_1899,FA_out_1899}=FA_cout_856+FA_out_869+FA_cout_917;
  assign {FA_cout_1900,FA_out_1900}=FA_out_858+FA_cout_884+FA_out_919;
  assign {FA_cout_1901,FA_out_1901}=FA_cout_859+FA_out_872+FA_cout_920;
  assign {FA_cout_1902,FA_out_1902}=FA_out_861+FA_cout_887+FA_out_922;
  assign {FA_cout_1903,FA_out_1903}=FA_cout_862+FA_out_875+FA_cout_923;
  assign {FA_cout_1904,FA_out_1904}=FA_out_864+FA_cout_890+FA_out_925;
  assign {FA_cout_1905,FA_out_1905}=FA_cout_865+FA_out_878+FA_cout_926;
  assign {FA_cout_1906,FA_out_1906}=FA_out_867+FA_cout_893+FA_out_928;
  assign {FA_cout_1907,FA_out_1907}=FA_cout_868+FA_out_881+FA_cout_929;
  assign {FA_cout_1908,FA_out_1908}=FA_out_835+HA_cout_14+FA_out_896;
  assign {FA_cout_1909,FA_out_1909}=FA_out_836+FA_cout_896+FA_out_897;
  assign {FA_cout_1910,FA_out_1910}=FA_out_837+FA_cout_897+FA_out_898;
  assign {FA_cout_1911,FA_out_1911}=FA_out_838+FA_cout_898+FA_out_899;
  assign {FA_cout_1912,FA_out_1912}=FA_out_839+FA_cout_899+FA_out_900;
  assign {FA_cout_1913,FA_out_1913}=FA_out_840+FA_cout_900+FA_out_901;
  assign {FA_cout_1914,FA_out_1914}=FA_out_841+FA_cout_901+FA_out_902;
  assign {FA_cout_1915,FA_out_1915}=FA_out_842+FA_cout_902+FA_out_903;
  assign {FA_cout_1916,FA_out_1916}=FA_out_843+FA_cout_903+FA_out_904;
  assign {FA_cout_1917,FA_out_1917}=FA_out_844+FA_cout_904+FA_out_905;
  assign {FA_cout_1918,FA_out_1918}=FA_out_845+FA_cout_905+FA_out_906;
  assign {FA_cout_1919,FA_out_1919}=FA_out_846+FA_cout_906+FA_out_907;
  assign {FA_cout_1920,FA_out_1920}=FA_out_847+FA_cout_907+FA_out_908;
  assign {FA_cout_1921,FA_out_1921}=FA_out_848+FA_cout_908+FA_out_909;
  assign {FA_cout_1922,FA_out_1922}=FA_out_849+FA_cout_909+FA_out_910;
  assign {FA_cout_1923,FA_out_1923}=FA_out_850+FA_cout_910+FA_out_911;
  assign {FA_cout_1924,FA_out_1924}=FA_out_851+FA_cout_911+FA_out_912;
  assign {FA_cout_1925,FA_out_1925}=FA_out_852+FA_cout_912+FA_out_913;
  assign {FA_cout_1926,FA_out_1926}=FA_out_853+FA_cout_913+FA_out_914;
  assign {FA_cout_1927,FA_out_1927}=FA_out_854+FA_cout_914+FA_out_915;
  assign {FA_cout_1928,FA_out_1928}=FA_out_855+FA_cout_915+FA_out_916;
  assign {FA_cout_1929,FA_out_1929}=FA_cout_869+FA_out_883+FA_cout_931;
  assign {FA_cout_1930,FA_out_1930}=FA_out_871+FA_cout_919+FA_out_933;
  assign {FA_cout_1931,FA_out_1931}=FA_cout_872+FA_out_886+FA_cout_934;
  assign {FA_cout_1932,FA_out_1932}=FA_out_874+FA_cout_922+FA_out_936;
  assign {FA_cout_1933,FA_out_1933}=FA_cout_875+FA_out_889+FA_cout_937;
  assign {FA_cout_1934,FA_out_1934}=FA_out_877+FA_cout_925+FA_out_939;
  assign {FA_cout_1935,FA_out_1935}=FA_cout_878+FA_out_892+FA_cout_940;
  assign {FA_cout_1936,FA_out_1936}=FA_out_880+FA_cout_928+FA_out_942;
  assign {FA_cout_1937,FA_out_1937}=FA_cout_881+FA_out_895+FA_cout_943;
  assign {FA_cout_1938,FA_out_1938}=FA_out_882+FA_cout_916+FA_out_945;
  assign {FA_cout_1939,FA_out_1939}=FA_cout_883+FA_out_918+FA_cout_946;
  assign {FA_cout_1940,FA_out_1940}=FA_out_885+FA_cout_933+FA_out_948;
  assign {FA_cout_1941,FA_out_1941}=FA_cout_886+FA_out_921+FA_cout_949;
  assign {FA_cout_1942,FA_out_1942}=FA_out_888+FA_cout_936+FA_out_951;
  assign {FA_cout_1943,FA_out_1943}=FA_cout_889+FA_out_924+FA_cout_952;
  assign {FA_cout_1944,FA_out_1944}=FA_out_891+FA_cout_939+FA_out_954;
  assign {FA_cout_1945,FA_out_1945}=FA_cout_892+FA_out_927+FA_cout_955;
  assign {FA_cout_1946,FA_out_1946}=FA_out_894+FA_cout_942+FA_out_957;
  assign {FA_cout_1947,FA_out_1947}=FA_cout_895+FA_out_930+FA_cout_958;
  assign {FA_cout_1948,FA_out_1948}=FA_out_917+FA_cout_945+FA_out_978;
  assign {FA_cout_1949,FA_out_1949}=FA_cout_918+FA_out_932+FA_cout_979;
  assign {FA_cout_1950,FA_out_1950}=FA_out_920+FA_cout_948+FA_out_981;
  assign {FA_cout_1951,FA_out_1951}=FA_cout_921+FA_out_935+FA_cout_982;
  assign {FA_cout_1952,FA_out_1952}=FA_out_923+FA_cout_951+FA_out_984;
  assign {FA_cout_1953,FA_out_1953}=FA_cout_924+FA_out_938+FA_cout_985;
  assign {FA_cout_1954,FA_out_1954}=FA_out_926+FA_cout_954+FA_out_987;
  assign {FA_cout_1955,FA_out_1955}=FA_cout_927+FA_out_941+FA_cout_988;
  assign {FA_cout_1956,FA_out_1956}=FA_out_929+FA_cout_957+FA_out_990;
  assign {FA_cout_1957,FA_out_1957}=FA_cout_930+FA_out_944+FA_cout_991;
  assign {FA_cout_1958,FA_out_1958}=FA_out_931+FA_cout_978+FA_out_993;
  assign {FA_cout_1959,FA_out_1959}=FA_cout_932+FA_out_947+FA_cout_994;
  assign {FA_cout_1960,FA_out_1960}=FA_out_934+FA_cout_981+FA_out_996;
  assign {FA_cout_1961,FA_out_1961}=FA_cout_935+FA_out_950+FA_cout_997;
  assign {FA_cout_1962,FA_out_1962}=FA_out_937+FA_cout_984+FA_out_999;
  assign {FA_cout_1963,FA_out_1963}=FA_cout_938+FA_out_953+FA_cout_1000;
  assign {FA_cout_1964,FA_out_1964}=FA_out_940+FA_cout_987+FA_out_1002;
  assign {FA_cout_1965,FA_out_1965}=FA_cout_941+FA_out_956+FA_cout_1003;
  assign {FA_cout_1966,FA_out_1966}=FA_out_943+FA_cout_990+FA_out_1005;
  assign {FA_cout_1967,FA_out_1967}=FA_cout_944+FA_out_959+FA_cout_1006;
  assign {FA_cout_1968,FA_out_1968}=FA_out_946+FA_cout_993+FA_out_1009;
  assign {FA_cout_1969,FA_out_1969}=FA_cout_947+FA_out_980+FA_cout_1010;
  assign {FA_cout_1970,FA_out_1970}=FA_out_949+FA_cout_996+FA_out_1012;
  assign {FA_cout_1971,FA_out_1971}=FA_cout_950+FA_out_983+FA_cout_1013;
  assign {FA_cout_1972,FA_out_1972}=FA_out_952+FA_cout_999+FA_out_1015;
  assign {FA_cout_1973,FA_out_1973}=FA_cout_953+FA_out_986+FA_cout_1016;
  assign {FA_cout_1974,FA_out_1974}=FA_out_955+FA_cout_1002+FA_out_1018;
  assign {FA_cout_1975,FA_out_1975}=FA_cout_956+FA_out_989+FA_cout_1019;
  assign {FA_cout_1976,FA_out_1976}=FA_out_958+FA_cout_1005+FA_out_1021;
  assign {FA_cout_1977,FA_out_1977}=FA_cout_959+FA_out_992+FA_cout_1022;
  assign {FA_cout_1978,FA_out_1978}=FA_cout_960+FA_out_961+inp_48[0];
  assign {FA_cout_1979,FA_out_1979}=FA_cout_961+FA_out_962+HA_out_16;
  assign {FA_cout_1980,FA_out_1980}=FA_cout_962+FA_out_963+HA_cout_16;
  assign {FA_cout_1981,FA_out_1981}=FA_cout_963+FA_out_964+FA_cout_1024;
  assign {FA_cout_1982,FA_out_1982}=FA_cout_964+FA_out_965+FA_cout_1025;
  assign {FA_cout_1983,FA_out_1983}=FA_cout_965+FA_out_966+FA_cout_1026;
  assign {FA_cout_1984,FA_out_1984}=FA_cout_966+FA_out_967+FA_cout_1027;
  assign {FA_cout_1985,FA_out_1985}=FA_cout_967+FA_out_968+FA_cout_1028;
  assign {FA_cout_1986,FA_out_1986}=FA_cout_968+FA_out_969+FA_cout_1029;
  assign {FA_cout_1987,FA_out_1987}=FA_cout_969+FA_out_970+FA_cout_1030;
  assign {FA_cout_1988,FA_out_1988}=FA_cout_970+FA_out_971+FA_cout_1031;
  assign {FA_cout_1989,FA_out_1989}=FA_cout_971+FA_out_972+FA_cout_1032;
  assign {FA_cout_1990,FA_out_1990}=FA_cout_972+FA_out_973+FA_cout_1033;
  assign {FA_cout_1991,FA_out_1991}=FA_cout_973+FA_out_974+FA_cout_1034;
  assign {FA_cout_1992,FA_out_1992}=FA_cout_974+FA_out_975+FA_cout_1035;
  assign {FA_cout_1993,FA_out_1993}=FA_cout_975+FA_out_976+FA_cout_1036;
  assign {FA_cout_1994,FA_out_1994}=FA_cout_976+FA_out_977+FA_cout_1037;
  assign {FA_cout_1995,FA_out_1995}=FA_cout_977+FA_out_1008+FA_cout_1038;
  assign {FA_cout_1996,FA_out_1996}=FA_out_979+FA_cout_1009+FA_out_1040;
  assign {FA_cout_1997,FA_out_1997}=FA_cout_980+FA_out_995+FA_cout_1041;
  assign {FA_cout_1998,FA_out_1998}=FA_out_982+FA_cout_1012+FA_out_1043;
  assign {FA_cout_1999,FA_out_1999}=FA_cout_983+FA_out_998+FA_cout_1044;
  assign {FA_cout_2000,FA_out_2000}=FA_out_985+FA_cout_1015+FA_out_1046;
  assign {FA_cout_2001,FA_out_2001}=FA_cout_986+FA_out_1001+FA_cout_1047;
  assign {FA_cout_2002,FA_out_2002}=FA_out_988+FA_cout_1018+FA_out_1049;
  assign {FA_cout_2003,FA_out_2003}=FA_cout_989+FA_out_1004+FA_cout_1050;
  assign {FA_cout_2004,FA_out_2004}=FA_out_991+FA_cout_1021+FA_out_1052;
  assign {FA_cout_2005,FA_out_2005}=FA_cout_992+FA_out_1007+FA_cout_1053;
  assign {FA_cout_2006,FA_out_2006}=FA_out_994+FA_cout_1040+FA_out_1056;
  assign {FA_cout_2007,FA_out_2007}=FA_cout_995+FA_out_1011+FA_cout_1057;
  assign {FA_cout_2008,FA_out_2008}=FA_out_997+FA_cout_1043+FA_out_1059;
  assign {FA_cout_2009,FA_out_2009}=FA_cout_998+FA_out_1014+FA_cout_1060;
  assign {FA_cout_2010,FA_out_2010}=FA_out_1000+FA_cout_1046+FA_out_1062;
  assign {FA_cout_2011,FA_out_2011}=FA_cout_1001+FA_out_1017+FA_cout_1063;
  assign {FA_cout_2012,FA_out_2012}=FA_out_1003+FA_cout_1049+FA_out_1065;
  assign {FA_cout_2013,FA_out_2013}=FA_cout_1004+FA_out_1020+FA_cout_1066;
  assign {FA_cout_2014,FA_out_2014}=FA_out_1006+FA_cout_1052+FA_out_1068;
  assign {FA_cout_2015,FA_out_2015}=FA_cout_1007+FA_out_1023+FA_cout_1069;
  assign {FA_cout_2016,FA_out_2016}=FA_cout_1008+FA_out_1039+FA_cout_1071;
  assign {FA_cout_2017,FA_out_2017}=FA_out_1010+FA_cout_1056+FA_out_1073;
  assign {FA_cout_2018,FA_out_2018}=FA_cout_1011+FA_out_1042+FA_cout_1074;
  assign {FA_cout_2019,FA_out_2019}=FA_out_1013+FA_cout_1059+FA_out_1076;
  assign {FA_cout_2020,FA_out_2020}=FA_cout_1014+FA_out_1045+FA_cout_1077;
  assign {FA_cout_2021,FA_out_2021}=FA_out_1016+FA_cout_1062+FA_out_1079;
  assign {FA_cout_2022,FA_out_2022}=FA_cout_1017+FA_out_1048+FA_cout_1080;
  assign {FA_cout_2023,FA_out_2023}=FA_out_1019+FA_cout_1065+FA_out_1082;
  assign {FA_cout_2024,FA_out_2024}=FA_cout_1020+FA_out_1051+FA_cout_1083;
  assign {FA_cout_2025,FA_out_2025}=FA_out_1022+FA_cout_1068+FA_out_1085;
  assign {FA_cout_2026,FA_out_2026}=FA_cout_1023+FA_out_1054+FA_cout_1086;
  assign {FA_cout_2027,FA_out_2027}=FA_cout_1039+FA_out_1055+FA_cout_1100;
  assign {FA_cout_2028,FA_out_2028}=FA_out_1041+FA_cout_1073+FA_out_1102;
  assign {FA_cout_2029,FA_out_2029}=FA_cout_1042+FA_out_1058+FA_cout_1103;
  assign {FA_cout_2030,FA_out_2030}=FA_out_1044+FA_cout_1076+FA_out_1105;
  assign {FA_cout_2031,FA_out_2031}=FA_cout_1045+FA_out_1061+FA_cout_1106;
  assign {FA_cout_2032,FA_out_2032}=FA_out_1047+FA_cout_1079+FA_out_1108;
  assign {FA_cout_2033,FA_out_2033}=FA_cout_1048+FA_out_1064+FA_cout_1109;
  assign {FA_cout_2034,FA_out_2034}=FA_out_1050+FA_cout_1082+FA_out_1111;
  assign {FA_cout_2035,FA_out_2035}=FA_cout_1051+FA_out_1067+FA_cout_1112;
  assign {FA_cout_2036,FA_out_2036}=FA_out_1053+FA_cout_1085+FA_out_1114;
  assign {FA_cout_2037,FA_out_2037}=FA_cout_1054+FA_out_1070+FA_cout_1115;
  assign {FA_cout_2038,FA_out_2038}=FA_out_1027+HA_cout_17+FA_out_1088;
  assign {FA_cout_2039,FA_out_2039}=FA_out_1028+FA_cout_1088+FA_out_1089;
  assign {FA_cout_2040,FA_out_2040}=FA_out_1029+FA_cout_1089+FA_out_1090;
  assign {FA_cout_2041,FA_out_2041}=FA_out_1030+FA_cout_1090+FA_out_1091;
  assign {FA_cout_2042,FA_out_2042}=FA_out_1031+FA_cout_1091+FA_out_1092;
  assign {FA_cout_2043,FA_out_2043}=FA_out_1032+FA_cout_1092+FA_out_1093;
  assign {FA_cout_2044,FA_out_2044}=FA_out_1033+FA_cout_1093+FA_out_1094;
  assign {FA_cout_2045,FA_out_2045}=FA_out_1034+FA_cout_1094+FA_out_1095;
  assign {FA_cout_2046,FA_out_2046}=FA_out_1035+FA_cout_1095+FA_out_1096;
  assign {FA_cout_2047,FA_out_2047}=FA_out_1036+FA_cout_1096+FA_out_1097;
  assign {FA_cout_2048,FA_out_2048}=FA_out_1037+FA_cout_1097+FA_out_1098;
  assign {FA_cout_2049,FA_out_2049}=FA_out_1038+FA_cout_1098+FA_out_1099;
  assign {FA_cout_2050,FA_out_2050}=FA_cout_1055+FA_out_1072+FA_cout_1117;
  assign {FA_cout_2051,FA_out_2051}=FA_out_1057+FA_cout_1102+FA_out_1119;
  assign {FA_cout_2052,FA_out_2052}=FA_cout_1058+FA_out_1075+FA_cout_1120;
  assign {FA_cout_2053,FA_out_2053}=FA_out_1060+FA_cout_1105+FA_out_1122;
  assign {FA_cout_2054,FA_out_2054}=FA_cout_1061+FA_out_1078+FA_cout_1123;
  assign {FA_cout_2055,FA_out_2055}=FA_out_1063+FA_cout_1108+FA_out_1125;
  assign {FA_cout_2056,FA_out_2056}=FA_cout_1064+FA_out_1081+FA_cout_1126;
  assign {FA_cout_2057,FA_out_2057}=FA_out_1066+FA_cout_1111+FA_out_1128;
  assign {FA_cout_2058,FA_out_2058}=FA_cout_1067+FA_out_1084+FA_cout_1129;
  assign {FA_cout_2059,FA_out_2059}=FA_out_1069+FA_cout_1114+FA_out_1131;
  assign {FA_cout_2060,FA_out_2060}=FA_cout_1070+FA_out_1087+FA_cout_1132;
  assign {FA_cout_2061,FA_out_2061}=FA_out_1071+FA_cout_1099+FA_out_1134;
  assign {FA_cout_2062,FA_out_2062}=FA_cout_1072+FA_out_1101+FA_cout_1135;
  assign {FA_cout_2063,FA_out_2063}=FA_out_1074+FA_cout_1119+FA_out_1137;
  assign {FA_cout_2064,FA_out_2064}=FA_cout_1075+FA_out_1104+FA_cout_1138;
  assign {FA_cout_2065,FA_out_2065}=FA_out_1077+FA_cout_1122+FA_out_1140;
  assign {FA_cout_2066,FA_out_2066}=FA_cout_1078+FA_out_1107+FA_cout_1141;
  assign {FA_cout_2067,FA_out_2067}=FA_out_1080+FA_cout_1125+FA_out_1143;
  assign {FA_cout_2068,FA_out_2068}=FA_cout_1081+FA_out_1110+FA_cout_1144;
  assign {FA_cout_2069,FA_out_2069}=FA_out_1083+FA_cout_1128+FA_out_1146;
  assign {FA_cout_2070,FA_out_2070}=FA_cout_1084+FA_out_1113+FA_cout_1147;
  assign {FA_cout_2071,FA_out_2071}=FA_out_1086+FA_cout_1131+FA_out_1149;
  assign {FA_cout_2072,FA_out_2072}=FA_cout_1087+FA_out_1116+FA_cout_1150;
  assign {FA_cout_2073,FA_out_2073}=FA_out_1100+FA_cout_1134+FA_out_1161;
  assign {FA_cout_2074,FA_out_2074}=FA_cout_1101+FA_out_1118+FA_cout_1162;
  assign {FA_cout_2075,FA_out_2075}=FA_out_1103+FA_cout_1137+FA_out_1164;
  assign {FA_cout_2076,FA_out_2076}=FA_cout_1104+FA_out_1121+FA_cout_1165;
  assign {FA_cout_2077,FA_out_2077}=FA_out_1106+FA_cout_1140+FA_out_1167;
  assign {FA_cout_2078,FA_out_2078}=FA_cout_1107+FA_out_1124+FA_cout_1168;
  assign {FA_cout_2079,FA_out_2079}=FA_out_1109+FA_cout_1143+FA_out_1170;
  assign {FA_cout_2080,FA_out_2080}=FA_cout_1110+FA_out_1127+FA_cout_1171;
  assign {FA_cout_2081,FA_out_2081}=FA_out_1112+FA_cout_1146+FA_out_1173;
  assign {FA_cout_2082,FA_out_2082}=FA_cout_1113+FA_out_1130+FA_cout_1174;
  assign {FA_cout_2083,FA_out_2083}=FA_out_1115+FA_cout_1149+FA_out_1176;
  assign {FA_cout_2084,FA_out_2084}=FA_cout_1116+FA_out_1133+FA_cout_1177;
  assign {FA_cout_2085,FA_out_2085}=FA_out_1117+FA_cout_1161+FA_out_1179;
  assign {FA_cout_2086,FA_out_2086}=FA_cout_1118+FA_out_1136+FA_cout_1180;
  assign {FA_cout_2087,FA_out_2087}=FA_out_1120+FA_cout_1164+FA_out_1182;
  assign {FA_cout_2088,FA_out_2088}=FA_cout_1121+FA_out_1139+FA_cout_1183;
  assign {FA_cout_2089,FA_out_2089}=FA_out_1123+FA_cout_1167+FA_out_1185;
  assign {FA_cout_2090,FA_out_2090}=FA_cout_1124+FA_out_1142+FA_cout_1186;
  assign {FA_cout_2091,FA_out_2091}=FA_out_1126+FA_cout_1170+FA_out_1188;
  assign {FA_cout_2092,FA_out_2092}=FA_cout_1127+FA_out_1145+FA_cout_1189;
  assign {FA_cout_2093,FA_out_2093}=FA_out_1129+FA_cout_1173+FA_out_1191;
  assign {FA_cout_2094,FA_out_2094}=FA_cout_1130+FA_out_1148+FA_cout_1192;
  assign {FA_cout_2095,FA_out_2095}=FA_out_1132+FA_cout_1176+FA_out_1194;
  assign {FA_cout_2096,FA_out_2096}=FA_cout_1133+FA_out_1151+FA_cout_1195;
  assign {FA_cout_2097,FA_out_2097}=FA_out_1135+FA_cout_1179+FA_out_1198;
  assign {FA_cout_2098,FA_out_2098}=FA_cout_1136+FA_out_1163+FA_cout_1199;
  assign {FA_cout_2099,FA_out_2099}=FA_out_1138+FA_cout_1182+FA_out_1201;
  assign {FA_cout_2100,FA_out_2100}=FA_cout_1139+FA_out_1166+FA_cout_1202;
  assign {FA_cout_2101,FA_out_2101}=FA_out_1141+FA_cout_1185+FA_out_1204;
  assign {FA_cout_2102,FA_out_2102}=FA_cout_1142+FA_out_1169+FA_cout_1205;
  assign {FA_cout_2103,FA_out_2103}=FA_out_1144+FA_cout_1188+FA_out_1207;
  assign {FA_cout_2104,FA_out_2104}=FA_cout_1145+FA_out_1172+FA_cout_1208;
  assign {FA_cout_2105,FA_out_2105}=FA_out_1147+FA_cout_1191+FA_out_1210;
  assign {FA_cout_2106,FA_out_2106}=FA_cout_1148+FA_out_1175+FA_cout_1211;
  assign {FA_cout_2107,FA_out_2107}=FA_out_1150+FA_cout_1194+FA_out_1213;
  assign {FA_cout_2108,FA_out_2108}=FA_cout_1151+FA_out_1178+FA_cout_1214;
  assign {FA_cout_2109,FA_out_2109}=FA_cout_1152+FA_out_1153+inp_57[0];
  assign {FA_cout_2110,FA_out_2110}=FA_cout_1153+FA_out_1154+HA_out_19;
  assign {FA_cout_2111,FA_out_2111}=FA_cout_1154+FA_out_1155+HA_cout_19;
  assign {FA_cout_2112,FA_out_2112}=FA_cout_1155+FA_out_1156+FA_cout_1216;
  assign {FA_cout_2113,FA_out_2113}=FA_cout_1156+FA_out_1157+FA_cout_1217;
  assign {FA_cout_2114,FA_out_2114}=FA_cout_1157+FA_out_1158+FA_cout_1218;
  assign {FA_cout_2115,FA_out_2115}=FA_cout_1158+FA_out_1159+FA_cout_1219;
  assign {FA_cout_2116,FA_out_2116}=FA_cout_1159+FA_out_1160+FA_cout_1220;
  assign {FA_cout_2117,FA_out_2117}=FA_cout_1160+FA_out_1197+FA_cout_1221;
  assign {FA_cout_2118,FA_out_2118}=FA_out_1162+FA_cout_1198+FA_out_1223;
  assign {FA_cout_2119,FA_out_2119}=FA_cout_1163+FA_out_1181+FA_cout_1224;
  assign {FA_cout_2120,FA_out_2120}=FA_out_1165+FA_cout_1201+FA_out_1226;
  assign {FA_cout_2121,FA_out_2121}=FA_cout_1166+FA_out_1184+FA_cout_1227;
  assign {FA_cout_2122,FA_out_2122}=FA_out_1168+FA_cout_1204+FA_out_1229;
  assign {FA_cout_2123,FA_out_2123}=FA_cout_1169+FA_out_1187+FA_cout_1230;
  assign {FA_cout_2124,FA_out_2124}=FA_out_1171+FA_cout_1207+FA_out_1232;
  assign {FA_cout_2125,FA_out_2125}=FA_cout_1172+FA_out_1190+FA_cout_1233;
  assign {FA_cout_2126,FA_out_2126}=FA_out_1174+FA_cout_1210+FA_out_1235;
  assign {FA_cout_2127,FA_out_2127}=FA_cout_1175+FA_out_1193+FA_cout_1236;
  assign {FA_cout_2128,FA_out_2128}=FA_out_1177+FA_cout_1213+FA_out_1238;
  assign {FA_cout_2129,FA_out_2129}=FA_cout_1178+FA_out_1196+FA_cout_1239;
  assign {FA_cout_2130,FA_out_2130}=FA_out_1180+FA_cout_1223+FA_out_1242;
  assign {FA_cout_2131,FA_out_2131}=FA_cout_1181+FA_out_1200+FA_cout_1243;
  assign {FA_cout_2132,FA_out_2132}=FA_out_1183+FA_cout_1226+FA_out_1245;
  assign {FA_cout_2133,FA_out_2133}=FA_cout_1184+FA_out_1203+FA_cout_1246;
  assign {FA_cout_2134,FA_out_2134}=FA_out_1186+FA_cout_1229+FA_out_1248;
  assign {FA_cout_2135,FA_out_2135}=FA_cout_1187+FA_out_1206+FA_cout_1249;
  assign {FA_cout_2136,FA_out_2136}=FA_out_1189+FA_cout_1232+FA_out_1251;
  assign {FA_cout_2137,FA_out_2137}=FA_cout_1190+FA_out_1209+FA_cout_1252;
  assign {FA_cout_2138,FA_out_2138}=FA_out_1192+FA_cout_1235+FA_out_1254;
  assign {FA_cout_2139,FA_out_2139}=FA_cout_1193+FA_out_1212+FA_cout_1255;
  assign {FA_cout_2140,FA_out_2140}=FA_out_1195+FA_cout_1238+FA_out_1257;
  assign {FA_cout_2141,FA_out_2141}=FA_cout_1196+FA_out_1215+FA_cout_1258;
  assign {FA_cout_2142,FA_out_2142}=FA_cout_1197+FA_out_1222+FA_cout_1260;
  assign {FA_cout_2143,FA_out_2143}=FA_out_1199+FA_cout_1242+FA_out_1262;
  assign {FA_cout_2144,FA_out_2144}=FA_cout_1200+FA_out_1225+FA_cout_1263;
  assign {FA_cout_2145,FA_out_2145}=FA_out_1202+FA_cout_1245+FA_out_1265;
  assign {FA_cout_2146,FA_out_2146}=FA_cout_1203+FA_out_1228+FA_cout_1266;
  assign {FA_cout_2147,FA_out_2147}=FA_out_1205+FA_cout_1248+FA_out_1268;
  assign {FA_cout_2148,FA_out_2148}=FA_cout_1206+FA_out_1231+FA_cout_1269;
  assign {FA_cout_2149,FA_out_2149}=FA_out_1208+FA_cout_1251+FA_out_1271;
  assign {FA_cout_2150,FA_out_2150}=FA_cout_1209+FA_out_1234+FA_cout_1272;
  assign {FA_cout_2151,FA_out_2151}=FA_out_1211+FA_cout_1254+FA_out_1274;
  assign {FA_cout_2152,FA_out_2152}=FA_cout_1212+FA_out_1237+FA_cout_1275;
  assign {FA_cout_2153,FA_out_2153}=FA_out_1214+FA_cout_1257+FA_out_1277;
  assign {FA_cout_2154,FA_out_2154}=FA_cout_1215+FA_out_1240+FA_cout_1278;
  assign {FA_cout_2155,FA_out_2155}=FA_cout_1222+FA_out_1241+FA_cout_1283;
  assign {FA_cout_2156,FA_out_2156}=FA_out_1224+FA_cout_1262+FA_out_1285;
  assign {FA_cout_2157,FA_out_2157}=FA_cout_1225+FA_out_1244+FA_cout_1286;
  assign {FA_cout_2158,FA_out_2158}=FA_out_1227+FA_cout_1265+FA_out_1288;
  assign {FA_cout_2159,FA_out_2159}=FA_cout_1228+FA_out_1247+FA_cout_1289;
  assign {FA_cout_2160,FA_out_2160}=FA_out_1230+FA_cout_1268+FA_out_1291;
  assign {FA_cout_2161,FA_out_2161}=FA_cout_1231+FA_out_1250+FA_cout_1292;
  assign {FA_cout_2162,FA_out_2162}=FA_out_1233+FA_cout_1271+FA_out_1294;
  assign {FA_cout_2163,FA_out_2163}=FA_cout_1234+FA_out_1253+FA_cout_1295;
  assign {FA_cout_2164,FA_out_2164}=FA_out_1236+FA_cout_1274+FA_out_1297;
  assign {FA_cout_2165,FA_out_2165}=FA_cout_1237+FA_out_1256+FA_cout_1298;
  assign {FA_cout_2166,FA_out_2166}=FA_out_1239+FA_cout_1277+FA_out_1300;
  assign {FA_cout_2167,FA_out_2167}=FA_cout_1240+FA_out_1259+FA_cout_1301;
  assign {FA_cout_2168,FA_out_2168}=FA_out_1219+HA_cout_20+FA_out_1280;
  assign {FA_cout_2169,FA_out_2169}=FA_out_1220+FA_cout_1280+FA_out_1281;
  assign {FA_cout_2170,FA_out_2170}=FA_out_1221+FA_cout_1281+FA_out_1282;
  assign {FA_cout_2171,FA_out_2171}=FA_cout_1241+FA_out_1261+FA_cout_1303;
  assign {FA_cout_2172,FA_out_2172}=FA_out_1243+FA_cout_1285+FA_out_1305;
  assign {FA_cout_2173,FA_out_2173}=FA_cout_1244+FA_out_1264+FA_cout_1306;
  assign {FA_cout_2174,FA_out_2174}=FA_out_1246+FA_cout_1288+FA_out_1308;
  assign {FA_cout_2175,FA_out_2175}=FA_cout_1247+FA_out_1267+FA_cout_1309;
  assign {FA_cout_2176,FA_out_2176}=FA_out_1249+FA_cout_1291+FA_out_1311;
  assign {FA_cout_2177,FA_out_2177}=FA_cout_1250+FA_out_1270+FA_cout_1312;
  assign {FA_cout_2178,FA_out_2178}=FA_out_1252+FA_cout_1294+FA_out_1314;
  assign {FA_cout_2179,FA_out_2179}=FA_cout_1253+FA_out_1273+FA_cout_1315;
  assign {FA_cout_2180,FA_out_2180}=FA_out_1255+FA_cout_1297+FA_out_1317;
  assign {FA_cout_2181,FA_out_2181}=FA_cout_1256+FA_out_1276+FA_cout_1318;
  assign {FA_cout_2182,FA_out_2182}=FA_out_1258+FA_cout_1300+FA_out_1320;
  assign {FA_cout_2183,FA_out_2183}=FA_cout_1259+FA_out_1279+FA_cout_1321;
  assign {FA_cout_2184,FA_out_2184}=FA_out_1260+FA_cout_1282+HA_out_21;
  assign {FA_cout_2185,FA_out_2185}=FA_cout_1261+FA_out_1284+HA_cout_22;
  assign {FA_cout_2186,FA_out_2186}=FA_out_1263+FA_cout_1305+HA_out_24;
  assign {FA_cout_2187,FA_out_2187}=FA_cout_1264+FA_out_1287+HA_cout_25;
  assign {FA_cout_2188,FA_out_2188}=FA_out_1266+FA_cout_1308+HA_out_27;
  assign {FA_cout_2189,FA_out_2189}=FA_cout_1267+FA_out_1290+HA_cout_28;
  assign {FA_cout_2190,FA_out_2190}=FA_out_1269+FA_cout_1311+HA_out_30;
  assign {FA_cout_2191,FA_out_2191}=FA_cout_1270+FA_out_1293+HA_cout_31;
  assign {FA_cout_2192,FA_out_2192}=FA_out_1272+FA_cout_1314+HA_out_33;
  assign {FA_cout_2193,FA_out_2193}=FA_cout_1273+FA_out_1296+HA_cout_34;
  assign {FA_cout_2194,FA_out_2194}=FA_out_1275+FA_cout_1317+HA_out_36;
  assign {FA_cout_2195,FA_out_2195}=FA_cout_1276+FA_out_1299+HA_cout_37;
  assign {FA_cout_2196,FA_out_2196}=FA_out_1278+FA_cout_1320+HA_out_39;
  assign {FA_cout_2197,FA_out_2197}=FA_cout_1279+FA_out_1302+HA_cout_40;
  assign {FA_cout_2198,FA_out_2198}=FA_out_1283+HA_cout_21+inp_63[3];
  assign {FA_cout_2199,FA_out_2199}=FA_out_1286+HA_cout_24+inp_63[12];
  assign {FA_cout_2200,FA_out_2200}=FA_out_1289+HA_cout_27+inp_63[21];
  assign {FA_cout_2201,FA_out_2201}=FA_out_1292+HA_cout_30+inp_63[30];
  assign {FA_cout_2202,FA_out_2202}=FA_out_1295+HA_cout_33+inp_63[39];
  assign {FA_cout_2203,FA_out_2203}=FA_out_1298+HA_cout_36+inp_63[48];
  assign {FA_cout_2204,FA_out_2204}=FA_out_1301+HA_cout_39+inp_63[57];
  assign {FA_cout_2205,FA_out_2205}=REGS_5+REGS_69+REGS_134;
  assign {FA_cout_2206,FA_out_2206}=REGS_6+REGS_70+REGS_135;
  assign {FA_cout_2207,FA_out_2207}=REGS_7+REGS_71+REGS_136;
  assign {FA_cout_2208,FA_out_2208}=REGS_8+REGS_72+REGS_137;
  assign {FA_cout_2209,FA_out_2209}=REGS_9+REGS_73+REGS_138;
  assign {FA_cout_2210,FA_out_2210}=REGS_10+REGS_74+REGS_139;
  assign {FA_cout_2211,FA_out_2211}=REGS_11+REGS_75+REGS_140;
  assign {FA_cout_2212,FA_out_2212}=REGS_12+REGS_76+REGS_141;
  assign {FA_cout_2213,FA_out_2213}=REGS_13+REGS_77+REGS_142;
  assign {FA_cout_2214,FA_out_2214}=REGS_14+REGS_78+REGS_143;
  assign {FA_cout_2215,FA_out_2215}=REGS_15+REGS_79+REGS_144;
  assign {FA_cout_2216,FA_out_2216}=REGS_16+REGS_80+REGS_145;
  assign {FA_cout_2217,FA_out_2217}=REGS_17+REGS_81+REGS_146;
  assign {FA_cout_2218,FA_out_2218}=REGS_18+REGS_82+REGS_147;
  assign {FA_cout_2219,FA_out_2219}=REGS_19+REGS_83+REGS_148;
  assign {FA_cout_2220,FA_out_2220}=REGS_20+REGS_84+REGS_149;
  assign {FA_cout_2221,FA_out_2221}=REGS_21+REGS_85+REGS_150;
  assign {FA_cout_2222,FA_out_2222}=REGS_22+REGS_86+REGS_151;
  assign {FA_cout_2223,FA_out_2223}=REGS_23+REGS_87+REGS_152;
  assign {FA_cout_2224,FA_out_2224}=REGS_24+REGS_88+REGS_153;
  assign {FA_cout_2225,FA_out_2225}=REGS_25+REGS_89+REGS_154;
  assign {FA_cout_2226,FA_out_2226}=REGS_26+REGS_90+REGS_155;
  assign {FA_cout_2227,FA_out_2227}=REGS_27+REGS_91+REGS_156;
  assign {FA_cout_2228,FA_out_2228}=REGS_28+REGS_92+REGS_157;
  assign {FA_cout_2229,FA_out_2229}=REGS_29+REGS_93+REGS_158;
  assign {FA_cout_2230,FA_out_2230}=REGS_30+REGS_94+REGS_159;
  assign {FA_cout_2231,FA_out_2231}=REGS_31+REGS_95+REGS_160;
  assign {FA_cout_2232,FA_out_2232}=REGS_32+REGS_96+REGS_161;
  assign {FA_cout_2233,FA_out_2233}=REGS_33+REGS_97+REGS_162;
  assign {FA_cout_2234,FA_out_2234}=REGS_34+REGS_98+REGS_163;
  assign {FA_cout_2235,FA_out_2235}=REGS_35+REGS_99+REGS_164;
  assign {FA_cout_2236,FA_out_2236}=REGS_36+REGS_100+REGS_165;
  assign {FA_cout_2237,FA_out_2237}=REGS_37+REGS_101+REGS_166;
  assign {FA_cout_2238,FA_out_2238}=REGS_38+REGS_102+REGS_167;
  assign {FA_cout_2239,FA_out_2239}=REGS_39+REGS_103+REGS_168;
  assign {FA_cout_2240,FA_out_2240}=REGS_40+REGS_104+REGS_169;
  assign {FA_cout_2241,FA_out_2241}=REGS_41+REGS_105+REGS_170;
  assign {FA_cout_2242,FA_out_2242}=REGS_42+REGS_106+REGS_171;
  assign {FA_cout_2243,FA_out_2243}=REGS_43+REGS_107+REGS_172;
  assign {FA_cout_2244,FA_out_2244}=REGS_44+REGS_108+REGS_173;
  assign {FA_cout_2245,FA_out_2245}=REGS_45+REGS_109+REGS_174;
  assign {FA_cout_2246,FA_out_2246}=REGS_46+REGS_110+REGS_175;
  assign {FA_cout_2247,FA_out_2247}=REGS_47+REGS_111+REGS_176;
  assign {FA_cout_2248,FA_out_2248}=REGS_48+REGS_112+REGS_177;
  assign {FA_cout_2249,FA_out_2249}=REGS_49+REGS_113+REGS_178;
  assign {FA_cout_2250,FA_out_2250}=REGS_50+REGS_114+REGS_179;
  assign {FA_cout_2251,FA_out_2251}=REGS_51+REGS_115+REGS_180;
  assign {FA_cout_2252,FA_out_2252}=REGS_52+REGS_116+REGS_181;
  assign {FA_cout_2253,FA_out_2253}=REGS_53+REGS_117+REGS_182;
  assign {FA_cout_2254,FA_out_2254}=REGS_54+REGS_118+REGS_183;
  assign {FA_cout_2255,FA_out_2255}=REGS_55+REGS_119+REGS_184;
  assign {FA_cout_2256,FA_out_2256}=REGS_56+REGS_120+REGS_185;
  assign {FA_cout_2257,FA_out_2257}=REGS_57+REGS_121+REGS_186;
  assign {FA_cout_2258,FA_out_2258}=REGS_58+REGS_122+REGS_187;
  assign {FA_cout_2259,FA_out_2259}=REGS_59+REGS_123+REGS_188;
  assign {FA_cout_2260,FA_out_2260}=REGS_60+REGS_124+REGS_189;
  assign {FA_cout_2261,FA_out_2261}=REGS_61+REGS_125+REGS_190;
  assign {FA_cout_2262,FA_out_2262}=REGS_62+REGS_126+REGS_191;
  assign {FA_cout_2263,FA_out_2263}=REGS_63+REGS_127+REGS_192;
  assign {FA_cout_2264,FA_out_2264}=REGS_64+REGS_128+REGS_193;
  assign {FA_cout_2265,FA_out_2265}=REGS_65+REGS_129+REGS_194;
  assign {FA_cout_2266,FA_out_2266}=REGS_66+REGS_130+REGS_256;
  assign {FA_cout_2267,FA_out_2267}=REGS_131+REGS_132+REGS_260;
  assign {FA_cout_2268,FA_out_2268}=REGS_133+REGS_195+REGS_264;
  assign {FA_cout_2269,FA_out_2269}=REGS_196+REGS_257+REGS_268;
  assign {FA_cout_2270,FA_out_2270}=REGS_202+REGS_274+REGS_333;
  assign {FA_cout_2271,FA_out_2271}=REGS_203+REGS_275+REGS_334;
  assign {FA_cout_2272,FA_out_2272}=REGS_204+REGS_276+REGS_335;
  assign {FA_cout_2273,FA_out_2273}=REGS_205+REGS_277+REGS_336;
  assign {FA_cout_2274,FA_out_2274}=REGS_206+REGS_278+REGS_337;
  assign {FA_cout_2275,FA_out_2275}=REGS_207+REGS_279+REGS_338;
  assign {FA_cout_2276,FA_out_2276}=REGS_208+REGS_280+REGS_339;
  assign {FA_cout_2277,FA_out_2277}=REGS_209+REGS_281+REGS_340;
  assign {FA_cout_2278,FA_out_2278}=REGS_210+REGS_282+REGS_341;
  assign {FA_cout_2279,FA_out_2279}=REGS_211+REGS_283+REGS_342;
  assign {FA_cout_2280,FA_out_2280}=REGS_212+REGS_284+REGS_343;
  assign {FA_cout_2281,FA_out_2281}=REGS_213+REGS_285+REGS_344;
  assign {FA_cout_2282,FA_out_2282}=REGS_214+REGS_286+REGS_345;
  assign {FA_cout_2283,FA_out_2283}=REGS_215+REGS_287+REGS_346;
  assign {FA_cout_2284,FA_out_2284}=REGS_216+REGS_288+REGS_347;
  assign {FA_cout_2285,FA_out_2285}=REGS_217+REGS_289+REGS_348;
  assign {FA_cout_2286,FA_out_2286}=REGS_218+REGS_290+REGS_349;
  assign {FA_cout_2287,FA_out_2287}=REGS_219+REGS_291+REGS_350;
  assign {FA_cout_2288,FA_out_2288}=REGS_220+REGS_292+REGS_351;
  assign {FA_cout_2289,FA_out_2289}=REGS_221+REGS_293+REGS_352;
  assign {FA_cout_2290,FA_out_2290}=REGS_222+REGS_294+REGS_353;
  assign {FA_cout_2291,FA_out_2291}=REGS_223+REGS_295+REGS_354;
  assign {FA_cout_2292,FA_out_2292}=REGS_224+REGS_296+REGS_355;
  assign {FA_cout_2293,FA_out_2293}=REGS_225+REGS_297+REGS_356;
  assign {FA_cout_2294,FA_out_2294}=REGS_226+REGS_298+REGS_357;
  assign {FA_cout_2295,FA_out_2295}=REGS_227+REGS_299+REGS_358;
  assign {FA_cout_2296,FA_out_2296}=REGS_228+REGS_300+REGS_359;
  assign {FA_cout_2297,FA_out_2297}=REGS_229+REGS_301+REGS_360;
  assign {FA_cout_2298,FA_out_2298}=REGS_230+REGS_302+REGS_361;
  assign {FA_cout_2299,FA_out_2299}=REGS_231+REGS_303+REGS_362;
  assign {FA_cout_2300,FA_out_2300}=REGS_232+REGS_304+REGS_363;
  assign {FA_cout_2301,FA_out_2301}=REGS_233+REGS_305+REGS_364;
  assign {FA_cout_2302,FA_out_2302}=REGS_234+REGS_306+REGS_365;
  assign {FA_cout_2303,FA_out_2303}=REGS_235+REGS_307+REGS_366;
  assign {FA_cout_2304,FA_out_2304}=REGS_236+REGS_308+REGS_367;
  assign {FA_cout_2305,FA_out_2305}=REGS_237+REGS_309+REGS_368;
  assign {FA_cout_2306,FA_out_2306}=REGS_238+REGS_310+REGS_369;
  assign {FA_cout_2307,FA_out_2307}=REGS_239+REGS_311+REGS_370;
  assign {FA_cout_2308,FA_out_2308}=REGS_240+REGS_312+REGS_371;
  assign {FA_cout_2309,FA_out_2309}=REGS_241+REGS_313+REGS_372;
  assign {FA_cout_2310,FA_out_2310}=REGS_242+REGS_314+REGS_373;
  assign {FA_cout_2311,FA_out_2311}=REGS_243+REGS_315+REGS_374;
  assign {FA_cout_2312,FA_out_2312}=REGS_244+REGS_316+REGS_375;
  assign {FA_cout_2313,FA_out_2313}=REGS_245+REGS_317+REGS_376;
  assign {FA_cout_2314,FA_out_2314}=REGS_246+REGS_318+REGS_377;
  assign {FA_cout_2315,FA_out_2315}=REGS_247+REGS_319+REGS_378;
  assign {FA_cout_2316,FA_out_2316}=REGS_248+REGS_320+REGS_379;
  assign {FA_cout_2317,FA_out_2317}=REGS_249+REGS_321+REGS_380;
  assign {FA_cout_2318,FA_out_2318}=REGS_250+REGS_322+REGS_381;
  assign {FA_cout_2319,FA_out_2319}=REGS_251+REGS_323+REGS_382;
  assign {FA_cout_2320,FA_out_2320}=REGS_252+REGS_324+REGS_383;
  assign {FA_cout_2321,FA_out_2321}=REGS_253+REGS_325+REGS_384;
  assign {FA_cout_2322,FA_out_2322}=REGS_254+REGS_326+REGS_385;
  assign {FA_cout_2323,FA_out_2323}=REGS_255+REGS_327+REGS_386;
  assign {FA_cout_2324,FA_out_2324}=REGS_258+REGS_261+REGS_330;
  assign {FA_cout_2325,FA_out_2325}=REGS_259+REGS_328+REGS_391;
  assign {FA_cout_2326,FA_out_2326}=REGS_262+REGS_265+REGS_388;
  assign {FA_cout_2327,FA_out_2327}=REGS_263+REGS_392+REGS_397;
  assign {FA_cout_2328,FA_out_2328}=REGS_266+REGS_269+REGS_394;
  assign {FA_cout_2329,FA_out_2329}=REGS_267+REGS_398+REGS_455;
  assign {FA_cout_2330,FA_out_2330}=REGS_270+REGS_331+REGS_400;
  assign {FA_cout_2331,FA_out_2331}=REGS_329+REGS_456+REGS_512;
  assign {FA_cout_2332,FA_out_2332}=REGS_332+REGS_389+REGS_458;
  assign {FA_cout_2333,FA_out_2333}=REGS_387+REGS_513+REGS_520;
  assign {FA_cout_2334,FA_out_2334}=REGS_390+REGS_395+REGS_515;
  assign {FA_cout_2335,FA_out_2335}=REGS_393+REGS_521+REGS_528;
  assign {FA_cout_2336,FA_out_2336}=REGS_396+REGS_401+REGS_523;
  assign {FA_cout_2337,FA_out_2337}=REGS_399+REGS_529+REGS_536;
  assign {FA_cout_2338,FA_out_2338}=REGS_402+REGS_459+REGS_531;
  assign {FA_cout_2339,FA_out_2339}=REGS_407+REGS_463+REGS_542;
  assign {FA_cout_2340,FA_out_2340}=REGS_408+REGS_464+REGS_543;
  assign {FA_cout_2341,FA_out_2341}=REGS_409+REGS_465+REGS_544;
  assign {FA_cout_2342,FA_out_2342}=REGS_410+REGS_466+REGS_545;
  assign {FA_cout_2343,FA_out_2343}=REGS_411+REGS_467+REGS_546;
  assign {FA_cout_2344,FA_out_2344}=REGS_412+REGS_468+REGS_547;
  assign {FA_cout_2345,FA_out_2345}=REGS_413+REGS_469+REGS_548;
  assign {FA_cout_2346,FA_out_2346}=REGS_414+REGS_470+REGS_549;
  assign {FA_cout_2347,FA_out_2347}=REGS_415+REGS_471+REGS_550;
  assign {FA_cout_2348,FA_out_2348}=REGS_416+REGS_472+REGS_551;
  assign {FA_cout_2349,FA_out_2349}=REGS_417+REGS_473+REGS_552;
  assign {FA_cout_2350,FA_out_2350}=REGS_418+REGS_474+REGS_553;
  assign {FA_cout_2351,FA_out_2351}=REGS_419+REGS_475+REGS_554;
  assign {FA_cout_2352,FA_out_2352}=REGS_420+REGS_476+REGS_555;
  assign {FA_cout_2353,FA_out_2353}=REGS_421+REGS_477+REGS_556;
  assign {FA_cout_2354,FA_out_2354}=REGS_422+REGS_478+REGS_557;
  assign {FA_cout_2355,FA_out_2355}=REGS_423+REGS_479+REGS_558;
  assign {FA_cout_2356,FA_out_2356}=REGS_424+REGS_480+REGS_559;
  assign {FA_cout_2357,FA_out_2357}=REGS_425+REGS_481+REGS_560;
  assign {FA_cout_2358,FA_out_2358}=REGS_426+REGS_482+REGS_561;
  assign {FA_cout_2359,FA_out_2359}=REGS_427+REGS_483+REGS_562;
  assign {FA_cout_2360,FA_out_2360}=REGS_428+REGS_484+REGS_563;
  assign {FA_cout_2361,FA_out_2361}=REGS_429+REGS_485+REGS_564;
  assign {FA_cout_2362,FA_out_2362}=REGS_430+REGS_486+REGS_565;
  assign {FA_cout_2363,FA_out_2363}=REGS_431+REGS_487+REGS_566;
  assign {FA_cout_2364,FA_out_2364}=REGS_432+REGS_488+REGS_567;
  assign {FA_cout_2365,FA_out_2365}=REGS_433+REGS_489+REGS_568;
  assign {FA_cout_2366,FA_out_2366}=REGS_434+REGS_490+REGS_569;
  assign {FA_cout_2367,FA_out_2367}=REGS_435+REGS_491+REGS_570;
  assign {FA_cout_2368,FA_out_2368}=REGS_436+REGS_492+REGS_571;
  assign {FA_cout_2369,FA_out_2369}=REGS_437+REGS_493+REGS_572;
  assign {FA_cout_2370,FA_out_2370}=REGS_438+REGS_494+REGS_573;
  assign {FA_cout_2371,FA_out_2371}=REGS_439+REGS_495+REGS_574;
  assign {FA_cout_2372,FA_out_2372}=REGS_440+REGS_496+REGS_575;
  assign {FA_cout_2373,FA_out_2373}=REGS_441+REGS_497+REGS_576;
  assign {FA_cout_2374,FA_out_2374}=REGS_442+REGS_498+REGS_577;
  assign {FA_cout_2375,FA_out_2375}=REGS_443+REGS_499+REGS_578;
  assign {FA_cout_2376,FA_out_2376}=REGS_444+REGS_500+REGS_579;
  assign {FA_cout_2377,FA_out_2377}=REGS_445+REGS_501+REGS_580;
  assign {FA_cout_2378,FA_out_2378}=REGS_446+REGS_502+REGS_581;
  assign {FA_cout_2379,FA_out_2379}=REGS_447+REGS_503+REGS_582;
  assign {FA_cout_2380,FA_out_2380}=REGS_448+REGS_504+REGS_583;
  assign {FA_cout_2381,FA_out_2381}=REGS_449+REGS_505+REGS_584;
  assign {FA_cout_2382,FA_out_2382}=REGS_450+REGS_506+REGS_585;
  assign {FA_cout_2383,FA_out_2383}=REGS_451+REGS_507+REGS_586;
  assign {FA_cout_2384,FA_out_2384}=REGS_452+REGS_508+REGS_587;
  assign {FA_cout_2385,FA_out_2385}=REGS_453+REGS_509+REGS_588;
  assign {FA_cout_2386,FA_out_2386}=REGS_454+REGS_510+REGS_589;
  assign {FA_cout_2387,FA_out_2387}=REGS_457+REGS_537+REGS_593;
  assign {FA_cout_2388,FA_out_2388}=REGS_460+REGS_516+REGS_539;
  assign {FA_cout_2389,FA_out_2389}=REGS_511+REGS_518+REGS_590;
  assign {FA_cout_2390,FA_out_2390}=REGS_514+REGS_594+REGS_646;
  assign {FA_cout_2391,FA_out_2391}=REGS_517+REGS_524+REGS_596;
  assign {FA_cout_2392,FA_out_2392}=REGS_519+REGS_526+REGS_653;
  assign {FA_cout_2393,FA_out_2393}=REGS_522+REGS_647+REGS_656;
  assign {FA_cout_2394,FA_out_2394}=REGS_525+REGS_532+REGS_649;
  assign {FA_cout_2395,FA_out_2395}=REGS_527+REGS_534+REGS_663;
  assign {FA_cout_2396,FA_out_2396}=REGS_530+REGS_657+REGS_666;
  assign {FA_cout_2397,FA_out_2397}=REGS_533+REGS_540+REGS_659;
  assign {FA_cout_2398,FA_out_2398}=REGS_535+REGS_591+REGS_716;
  assign {FA_cout_2399,FA_out_2399}=REGS_538+REGS_667+REGS_719;
  assign {FA_cout_2400,FA_out_2400}=REGS_541+REGS_597+REGS_669;
  assign {FA_cout_2401,FA_out_2401}=REGS_592+REGS_644+REGS_768;
  assign {FA_cout_2402,FA_out_2402}=REGS_595+REGS_720+REGS_771;
  assign {FA_cout_2403,FA_out_2403}=REGS_598+REGS_650+REGS_722;
  assign {FA_cout_2404,FA_out_2404}=REGS_603+REGS_674+REGS_725;
  assign {FA_cout_2405,FA_out_2405}=REGS_604+REGS_675+REGS_726;
  assign {FA_cout_2406,FA_out_2406}=REGS_605+REGS_676+REGS_727;
  assign {FA_cout_2407,FA_out_2407}=REGS_606+REGS_677+REGS_728;
  assign {FA_cout_2408,FA_out_2408}=REGS_607+REGS_678+REGS_729;
  assign {FA_cout_2409,FA_out_2409}=REGS_608+REGS_679+REGS_730;
  assign {FA_cout_2410,FA_out_2410}=REGS_609+REGS_680+REGS_731;
  assign {FA_cout_2411,FA_out_2411}=REGS_610+REGS_681+REGS_732;
  assign {FA_cout_2412,FA_out_2412}=REGS_611+REGS_682+REGS_733;
  assign {FA_cout_2413,FA_out_2413}=REGS_612+REGS_683+REGS_734;
  assign {FA_cout_2414,FA_out_2414}=REGS_613+REGS_684+REGS_735;
  assign {FA_cout_2415,FA_out_2415}=REGS_614+REGS_685+REGS_736;
  assign {FA_cout_2416,FA_out_2416}=REGS_615+REGS_686+REGS_737;
  assign {FA_cout_2417,FA_out_2417}=REGS_616+REGS_687+REGS_738;
  assign {FA_cout_2418,FA_out_2418}=REGS_617+REGS_688+REGS_739;
  assign {FA_cout_2419,FA_out_2419}=REGS_618+REGS_689+REGS_740;
  assign {FA_cout_2420,FA_out_2420}=REGS_619+REGS_690+REGS_741;
  assign {FA_cout_2421,FA_out_2421}=REGS_620+REGS_691+REGS_742;
  assign {FA_cout_2422,FA_out_2422}=REGS_621+REGS_692+REGS_743;
  assign {FA_cout_2423,FA_out_2423}=REGS_622+REGS_693+REGS_744;
  assign {FA_cout_2424,FA_out_2424}=REGS_623+REGS_694+REGS_745;
  assign {FA_cout_2425,FA_out_2425}=REGS_624+REGS_695+REGS_746;
  assign {FA_cout_2426,FA_out_2426}=REGS_625+REGS_696+REGS_747;
  assign {FA_cout_2427,FA_out_2427}=REGS_626+REGS_697+REGS_748;
  assign {FA_cout_2428,FA_out_2428}=REGS_627+REGS_698+REGS_749;
  assign {FA_cout_2429,FA_out_2429}=REGS_628+REGS_699+REGS_750;
  assign {FA_cout_2430,FA_out_2430}=REGS_629+REGS_700+REGS_751;
  assign {FA_cout_2431,FA_out_2431}=REGS_630+REGS_701+REGS_752;
  assign {FA_cout_2432,FA_out_2432}=REGS_631+REGS_702+REGS_753;
  assign {FA_cout_2433,FA_out_2433}=REGS_632+REGS_703+REGS_754;
  assign {FA_cout_2434,FA_out_2434}=REGS_633+REGS_704+REGS_755;
  assign {FA_cout_2435,FA_out_2435}=REGS_634+REGS_705+REGS_756;
  assign {FA_cout_2436,FA_out_2436}=REGS_635+REGS_706+REGS_757;
  assign {FA_cout_2437,FA_out_2437}=REGS_636+REGS_707+REGS_758;
  assign {FA_cout_2438,FA_out_2438}=REGS_637+REGS_708+REGS_759;
  assign {FA_cout_2439,FA_out_2439}=REGS_638+REGS_709+REGS_760;
  assign {FA_cout_2440,FA_out_2440}=REGS_639+REGS_710+REGS_761;
  assign {FA_cout_2441,FA_out_2441}=REGS_640+REGS_711+REGS_762;
  assign {FA_cout_2442,FA_out_2442}=REGS_641+REGS_712+REGS_763;
  assign {FA_cout_2443,FA_out_2443}=REGS_642+REGS_713+REGS_764;
  assign {FA_cout_2444,FA_out_2444}=REGS_643+REGS_714+REGS_765;
  assign {FA_cout_2445,FA_out_2445}=REGS_645+REGS_654+REGS_780;
  assign {FA_cout_2446,FA_out_2446}=REGS_648+REGS_772+REGS_783;
  assign {FA_cout_2447,FA_out_2447}=REGS_651+REGS_660+REGS_774;
  assign {FA_cout_2448,FA_out_2448}=REGS_652+REGS_766+REGS_777;
  assign {FA_cout_2449,FA_out_2449}=REGS_655+REGS_664+REGS_792;
  assign {FA_cout_2450,FA_out_2450}=REGS_658+REGS_784+REGS_795;
  assign {FA_cout_2451,FA_out_2451}=REGS_661+REGS_670+REGS_786;
  assign {FA_cout_2452,FA_out_2452}=REGS_662+REGS_778+REGS_789;
  assign {FA_cout_2453,FA_out_2453}=REGS_665+REGS_717+REGS_804;
  assign {FA_cout_2454,FA_out_2454}=REGS_668+REGS_796+REGS_807;
  assign {FA_cout_2455,FA_out_2455}=REGS_671+REGS_723+REGS_798;
  assign {FA_cout_2456,FA_out_2456}=REGS_715+REGS_790+REGS_801;
  assign {FA_cout_2457,FA_out_2457}=REGS_718+REGS_769+REGS_856;
  assign {FA_cout_2458,FA_out_2458}=REGS_721+REGS_808+REGS_859;
  assign {FA_cout_2459,FA_out_2459}=REGS_724+REGS_775+REGS_810;
  assign {FA_cout_2460,FA_out_2460}=REGS_767+REGS_802+REGS_853;
  assign {FA_cout_2461,FA_out_2461}=REGS_770+REGS_781+REGS_904;
  assign {FA_cout_2462,FA_out_2462}=REGS_773+REGS_860+REGS_907;
  assign {FA_cout_2463,FA_out_2463}=REGS_776+REGS_787+REGS_862;
  assign {FA_cout_2464,FA_out_2464}=REGS_779+REGS_854+REGS_901;
  assign {FA_cout_2465,FA_out_2465}=REGS_782+REGS_793+REGS_918;
  assign {FA_cout_2466,FA_out_2466}=REGS_785+REGS_908+REGS_921;
  assign {FA_cout_2467,FA_out_2467}=REGS_788+REGS_799+REGS_910;
  assign {FA_cout_2468,FA_out_2468}=REGS_791+REGS_902+REGS_915;
  assign {FA_cout_2469,FA_out_2469}=REGS_794+REGS_805+REGS_932;
  assign {FA_cout_2470,FA_out_2470}=REGS_797+REGS_922+REGS_935;
  assign {FA_cout_2471,FA_out_2471}=REGS_800+REGS_811+REGS_924;
  assign {FA_cout_2472,FA_out_2472}=REGS_803+REGS_916+REGS_929;
  assign {FA_cout_2473,FA_out_2473}=REGS_806+REGS_857+REGS_980;
  assign {FA_cout_2474,FA_out_2474}=REGS_809+REGS_936+REGS_983;
  assign {FA_cout_2475,FA_out_2475}=REGS_812+REGS_863+REGS_938;
  assign {FA_cout_2476,FA_out_2476}=REGS_818+REGS_867+REGS_941;
  assign {FA_cout_2477,FA_out_2477}=REGS_819+REGS_868+REGS_942;
  assign {FA_cout_2478,FA_out_2478}=REGS_820+REGS_869+REGS_943;
  assign {FA_cout_2479,FA_out_2479}=REGS_821+REGS_870+REGS_944;
  assign {FA_cout_2480,FA_out_2480}=REGS_822+REGS_871+REGS_945;
  assign {FA_cout_2481,FA_out_2481}=REGS_823+REGS_872+REGS_946;
  assign {FA_cout_2482,FA_out_2482}=REGS_824+REGS_873+REGS_947;
  assign {FA_cout_2483,FA_out_2483}=REGS_825+REGS_874+REGS_948;
  assign {FA_cout_2484,FA_out_2484}=REGS_826+REGS_875+REGS_949;
  assign {FA_cout_2485,FA_out_2485}=REGS_827+REGS_876+REGS_950;
  assign {FA_cout_2486,FA_out_2486}=REGS_828+REGS_877+REGS_951;
  assign {FA_cout_2487,FA_out_2487}=REGS_829+REGS_878+REGS_952;
  assign {FA_cout_2488,FA_out_2488}=REGS_830+REGS_879+REGS_953;
  assign {FA_cout_2489,FA_out_2489}=REGS_831+REGS_880+REGS_954;
  assign {FA_cout_2490,FA_out_2490}=REGS_832+REGS_881+REGS_955;
  assign {FA_cout_2491,FA_out_2491}=REGS_833+REGS_882+REGS_956;
  assign {FA_cout_2492,FA_out_2492}=REGS_834+REGS_883+REGS_957;
  assign {FA_cout_2493,FA_out_2493}=REGS_835+REGS_884+REGS_958;
  assign {FA_cout_2494,FA_out_2494}=REGS_836+REGS_885+REGS_959;
  assign {FA_cout_2495,FA_out_2495}=REGS_837+REGS_886+REGS_960;
  assign {FA_cout_2496,FA_out_2496}=REGS_838+REGS_887+REGS_961;
  assign {FA_cout_2497,FA_out_2497}=REGS_839+REGS_888+REGS_962;
  assign {FA_cout_2498,FA_out_2498}=REGS_840+REGS_889+REGS_963;
  assign {FA_cout_2499,FA_out_2499}=REGS_841+REGS_890+REGS_964;
  assign {FA_cout_2500,FA_out_2500}=REGS_842+REGS_891+REGS_965;
  assign {FA_cout_2501,FA_out_2501}=REGS_843+REGS_892+REGS_966;
  assign {FA_cout_2502,FA_out_2502}=REGS_844+REGS_893+REGS_967;
  assign {FA_cout_2503,FA_out_2503}=REGS_845+REGS_894+REGS_968;
  assign {FA_cout_2504,FA_out_2504}=REGS_846+REGS_895+REGS_969;
  assign {FA_cout_2505,FA_out_2505}=REGS_847+REGS_896+REGS_970;
  assign {FA_cout_2506,FA_out_2506}=REGS_848+REGS_897+REGS_971;
  assign {FA_cout_2507,FA_out_2507}=REGS_849+REGS_898+REGS_972;
  assign {FA_cout_2508,FA_out_2508}=REGS_850+REGS_899+REGS_973;
  assign {FA_cout_2509,FA_out_2509}=REGS_851+REGS_900+REGS_974;
  assign {FA_cout_2510,FA_out_2510}=REGS_852+REGS_913+REGS_1022;
  assign {FA_cout_2511,FA_out_2511}=REGS_855+REGS_930+REGS_977;
  assign {FA_cout_2512,FA_out_2512}=REGS_858+REGS_905+REGS_1028;
  assign {FA_cout_2513,FA_out_2513}=REGS_861+REGS_984+REGS_1031;
  assign {FA_cout_2514,FA_out_2514}=REGS_864+REGS_911+REGS_986;
  assign {FA_cout_2515,FA_out_2515}=REGS_903+REGS_978+REGS_1025;
  assign {FA_cout_2516,FA_out_2516}=REGS_906+REGS_919+REGS_1044;
  assign {FA_cout_2517,FA_out_2517}=REGS_909+REGS_1032+REGS_1047;
  assign {FA_cout_2518,FA_out_2518}=REGS_912+REGS_925+REGS_1034;
  assign {FA_cout_2519,FA_out_2519}=REGS_914+REGS_927+REGS_1038;
  assign {FA_cout_2520,FA_out_2520}=REGS_917+REGS_1026+REGS_1041;
  assign {FA_cout_2521,FA_out_2521}=REGS_920+REGS_933+REGS_1060;
  assign {FA_cout_2522,FA_out_2522}=REGS_923+REGS_1048+REGS_1063;
  assign {FA_cout_2523,FA_out_2523}=REGS_926+REGS_939+REGS_1050;
  assign {FA_cout_2524,FA_out_2524}=REGS_928+REGS_975+REGS_1054;
  assign {FA_cout_2525,FA_out_2525}=REGS_931+REGS_1042+REGS_1057;
  assign {FA_cout_2526,FA_out_2526}=REGS_934+REGS_981+REGS_1076;
  assign {FA_cout_2527,FA_out_2527}=REGS_937+REGS_1064+REGS_1079;
  assign {FA_cout_2528,FA_out_2528}=REGS_940+REGS_987+REGS_1066;
  assign {FA_cout_2529,FA_out_2529}=REGS_976+REGS_1023+REGS_1070;
  assign {FA_cout_2530,FA_out_2530}=REGS_979+REGS_1058+REGS_1073;
  assign {FA_cout_2531,FA_out_2531}=REGS_982+REGS_1029+REGS_1123;
  assign {FA_cout_2532,FA_out_2532}=REGS_985+REGS_1080+REGS_1126;
  assign {FA_cout_2533,FA_out_2533}=REGS_988+REGS_1035+REGS_1082;
  assign {FA_cout_2534,FA_out_2534}=REGS_995+REGS_1088+REGS_1132;
  assign {FA_cout_2535,FA_out_2535}=REGS_996+REGS_1089+REGS_1133;
  assign {FA_cout_2536,FA_out_2536}=REGS_997+REGS_1090+REGS_1134;
  assign {FA_cout_2537,FA_out_2537}=REGS_998+REGS_1091+REGS_1135;
  assign {FA_cout_2538,FA_out_2538}=REGS_999+REGS_1092+REGS_1136;
  assign {FA_cout_2539,FA_out_2539}=REGS_1000+REGS_1093+REGS_1137;
  assign {FA_cout_2540,FA_out_2540}=REGS_1001+REGS_1094+REGS_1138;
  assign {FA_cout_2541,FA_out_2541}=REGS_1002+REGS_1095+REGS_1139;
  assign {FA_cout_2542,FA_out_2542}=REGS_1003+REGS_1096+REGS_1140;
  assign {FA_cout_2543,FA_out_2543}=REGS_1004+REGS_1097+REGS_1141;
  assign {FA_cout_2544,FA_out_2544}=REGS_1005+REGS_1098+REGS_1142;
  assign {FA_cout_2545,FA_out_2545}=REGS_1006+REGS_1099+REGS_1143;
  assign {FA_cout_2546,FA_out_2546}=REGS_1007+REGS_1100+REGS_1144;
  assign {FA_cout_2547,FA_out_2547}=REGS_1008+REGS_1101+REGS_1145;
  assign {FA_cout_2548,FA_out_2548}=REGS_1009+REGS_1102+REGS_1146;
  assign {FA_cout_2549,FA_out_2549}=REGS_1010+REGS_1103+REGS_1147;
  assign {FA_cout_2550,FA_out_2550}=REGS_1011+REGS_1104+REGS_1148;
  assign {FA_cout_2551,FA_out_2551}=REGS_1012+REGS_1105+REGS_1149;
  assign {FA_cout_2552,FA_out_2552}=REGS_1013+REGS_1106+REGS_1150;
  assign {FA_cout_2553,FA_out_2553}=REGS_1014+REGS_1107+REGS_1151;
  assign {FA_cout_2554,FA_out_2554}=REGS_1015+REGS_1108+REGS_1152;
  assign {FA_cout_2555,FA_out_2555}=REGS_1016+REGS_1109+REGS_1153;
  assign {FA_cout_2556,FA_out_2556}=REGS_1017+REGS_1110+REGS_1154;
  assign {FA_cout_2557,FA_out_2557}=REGS_1018+REGS_1111+REGS_1155;
  assign {FA_cout_2558,FA_out_2558}=REGS_1019+REGS_1112+REGS_1156;
  assign {FA_cout_2559,FA_out_2559}=REGS_1020+REGS_1113+REGS_1157;
  assign {FA_cout_2560,FA_out_2560}=REGS_1021+REGS_1114+REGS_1158;
  assign {FA_cout_2561,FA_out_2561}=REGS_1024+REGS_1039+REGS_1117;
  assign {FA_cout_2562,FA_out_2562}=REGS_1027+REGS_1074+REGS_1120;
  assign {FA_cout_2563,FA_out_2563}=REGS_1030+REGS_1045+REGS_1166;
  assign {FA_cout_2564,FA_out_2564}=REGS_1033+REGS_1127+REGS_1169;
  assign {FA_cout_2565,FA_out_2565}=REGS_1036+REGS_1051+REGS_1129;
  assign {FA_cout_2566,FA_out_2566}=REGS_1037+REGS_1115+REGS_1175;
  assign {FA_cout_2567,FA_out_2567}=REGS_1040+REGS_1055+REGS_1160;
  assign {FA_cout_2568,FA_out_2568}=REGS_1043+REGS_1121+REGS_1163;
  assign {FA_cout_2569,FA_out_2569}=REGS_1046+REGS_1061+REGS_1184;
  assign {FA_cout_2570,FA_out_2570}=REGS_1049+REGS_1170+REGS_1187;
  assign {FA_cout_2571,FA_out_2571}=REGS_1052+REGS_1067+REGS_1172;
  assign {FA_cout_2572,FA_out_2572}=REGS_1053+REGS_1176+REGS_1193;
  assign {FA_cout_2573,FA_out_2573}=REGS_1056+REGS_1071+REGS_1178;
  assign {FA_cout_2574,FA_out_2574}=REGS_1059+REGS_1164+REGS_1181;
  assign {FA_cout_2575,FA_out_2575}=REGS_1062+REGS_1077+REGS_1202;
  assign {FA_cout_2576,FA_out_2576}=REGS_1065+REGS_1188+REGS_1205;
  assign {FA_cout_2577,FA_out_2577}=REGS_1068+REGS_1083+REGS_1190;
  assign {FA_cout_2578,FA_out_2578}=REGS_1069+REGS_1194+REGS_1236;
  assign {FA_cout_2579,FA_out_2579}=REGS_1072+REGS_1118+REGS_1196;
  assign {FA_cout_2580,FA_out_2580}=REGS_1075+REGS_1182+REGS_1199;
  assign {FA_cout_2581,FA_out_2581}=REGS_1078+REGS_1124+REGS_1245;
  assign {FA_cout_2582,FA_out_2582}=REGS_1081+REGS_1206+REGS_1248;
  assign {FA_cout_2583,FA_out_2583}=REGS_1084+REGS_1130+REGS_1208;
  assign {FA_cout_2584,FA_out_2584}=REGS_1116+REGS_1237+REGS_1278;
  assign {FA_cout_2585,FA_out_2585}=REGS_1119+REGS_1161+REGS_1239;
  assign {FA_cout_2586,FA_out_2586}=REGS_1122+REGS_1200+REGS_1242;
  assign {FA_cout_2587,FA_out_2587}=REGS_1125+REGS_1167+REGS_1287;
  assign {FA_cout_2588,FA_out_2588}=REGS_1128+REGS_1249+REGS_1290;
  assign {FA_cout_2589,FA_out_2589}=REGS_1131+REGS_1173+REGS_1251;
  assign {FA_cout_2590,FA_out_2590}=REGS_1159+REGS_1279+REGS_1298;
  assign {FA_cout_2591,FA_out_2591}=REGS_1162+REGS_1179+REGS_1281;
  assign {FA_cout_2592,FA_out_2592}=REGS_1165+REGS_1243+REGS_1284;
  assign {FA_cout_2593,FA_out_2593}=REGS_1168+REGS_1185+REGS_1307;
  assign {FA_cout_2594,FA_out_2594}=REGS_1171+REGS_1291+REGS_1310;
  assign {FA_cout_2595,FA_out_2595}=REGS_1174+REGS_1191+REGS_1293;
  assign {FA_cout_2596,FA_out_2596}=REGS_1177+REGS_1299+REGS_1318;
  assign {FA_cout_2597,FA_out_2597}=REGS_1180+REGS_1197+REGS_1301;
  assign {FA_cout_2598,FA_out_2598}=REGS_1183+REGS_1285+REGS_1304;
  assign {FA_cout_2599,FA_out_2599}=REGS_1186+REGS_1203+REGS_1327;
  assign {FA_cout_2600,FA_out_2600}=REGS_1189+REGS_1311+REGS_1330;
  assign {FA_cout_2601,FA_out_2601}=REGS_1192+REGS_1209+REGS_1313;
  assign {FA_cout_2602,FA_out_2602}=REGS_1195+REGS_1319+REGS_1338;
  assign {FA_cout_2603,FA_out_2603}=REGS_1198+REGS_1240+REGS_1321;
  assign {FA_cout_2604,FA_out_2604}=REGS_1201+REGS_1305+REGS_1324;
  assign {FA_cout_2605,FA_out_2605}=REGS_1204+REGS_1246+REGS_1347;
  assign {FA_cout_2606,FA_out_2606}=REGS_1207+REGS_1331+REGS_1350;
  assign {FA_cout_2607,FA_out_2607}=REGS_1210+REGS_1252+REGS_1333;
  assign {FA_cout_2608,FA_out_2608}=REGS_1215+REGS_1256+REGS_1356;
  assign {FA_cout_2609,FA_out_2609}=REGS_1216+REGS_1257+REGS_1357;
  assign {FA_cout_2610,FA_out_2610}=REGS_1217+REGS_1258+REGS_1358;
  assign {FA_cout_2611,FA_out_2611}=REGS_1218+REGS_1259+REGS_1359;
  assign {FA_cout_2612,FA_out_2612}=REGS_1219+REGS_1260+REGS_1360;
  assign {FA_cout_2613,FA_out_2613}=REGS_1220+REGS_1261+REGS_1361;
  assign {FA_cout_2614,FA_out_2614}=REGS_1221+REGS_1262+REGS_1362;
  assign {FA_cout_2615,FA_out_2615}=REGS_1222+REGS_1263+REGS_1363;
  assign {FA_cout_2616,FA_out_2616}=REGS_1223+REGS_1264+REGS_1364;
  assign {FA_cout_2617,FA_out_2617}=REGS_1224+REGS_1265+REGS_1365;
  assign {FA_cout_2618,FA_out_2618}=REGS_1225+REGS_1266+REGS_1366;
  assign {FA_cout_2619,FA_out_2619}=REGS_1226+REGS_1267+REGS_1367;
  assign {FA_cout_2620,FA_out_2620}=REGS_1227+REGS_1268+REGS_1368;
  assign {FA_cout_2621,FA_out_2621}=REGS_1228+REGS_1269+REGS_1369;
  assign {FA_cout_2622,FA_out_2622}=REGS_1229+REGS_1270+REGS_1370;
  assign {FA_cout_2623,FA_out_2623}=REGS_1230+REGS_1271+REGS_1371;
  assign {FA_cout_2624,FA_out_2624}=REGS_1231+REGS_1272+REGS_1372;
  assign {FA_cout_2625,FA_out_2625}=REGS_1232+REGS_1273+REGS_1373;
  assign {FA_cout_2626,FA_out_2626}=REGS_1233+REGS_1274+REGS_1374;
  assign {FA_cout_2627,FA_out_2627}=REGS_1234+REGS_1275+REGS_1375;
  assign {FA_cout_2628,FA_out_2628}=REGS_1235+REGS_1276+REGS_1376;
  assign {FA_cout_2629,FA_out_2629}=REGS_1238+REGS_1339+REGS_1380;
  assign {FA_cout_2630,FA_out_2630}=REGS_1241+REGS_1282+REGS_1341;
  assign {FA_cout_2631,FA_out_2631}=REGS_1244+REGS_1325+REGS_1344;
  assign {FA_cout_2632,FA_out_2632}=REGS_1247+REGS_1288+REGS_1389;
  assign {FA_cout_2633,FA_out_2633}=REGS_1250+REGS_1351+REGS_1392;
  assign {FA_cout_2634,FA_out_2634}=REGS_1253+REGS_1294+REGS_1353;
  assign {FA_cout_2635,FA_out_2635}=REGS_1277+REGS_1296+REGS_1377;
  assign {FA_cout_2636,FA_out_2636}=REGS_1280+REGS_1381+REGS_1418;
  assign {FA_cout_2637,FA_out_2637}=REGS_1283+REGS_1302+REGS_1383;
  assign {FA_cout_2638,FA_out_2638}=REGS_1286+REGS_1345+REGS_1386;
  assign {FA_cout_2639,FA_out_2639}=REGS_1289+REGS_1308+REGS_1427;
  assign {FA_cout_2640,FA_out_2640}=REGS_1292+REGS_1393+REGS_1430;
  assign {FA_cout_2641,FA_out_2641}=REGS_1295+REGS_1314+REGS_1395;
  assign {FA_cout_2642,FA_out_2642}=REGS_1297+REGS_1316+REGS_1437;
  assign {FA_cout_2643,FA_out_2643}=REGS_1300+REGS_1419+REGS_1440;
  assign {FA_cout_2644,FA_out_2644}=REGS_1303+REGS_1322+REGS_1421;
  assign {FA_cout_2645,FA_out_2645}=REGS_1306+REGS_1387+REGS_1424;
  assign {FA_cout_2646,FA_out_2646}=REGS_1309+REGS_1328+REGS_1449;
  assign {FA_cout_2647,FA_out_2647}=REGS_1312+REGS_1431+REGS_1452;
  assign {FA_cout_2648,FA_out_2648}=REGS_1315+REGS_1334+REGS_1433;
  assign {FA_cout_2649,FA_out_2649}=REGS_1317+REGS_1336+REGS_1459;
  assign {FA_cout_2650,FA_out_2650}=REGS_1320+REGS_1441+REGS_1462;
  assign {FA_cout_2651,FA_out_2651}=REGS_1323+REGS_1342+REGS_1443;
  assign {FA_cout_2652,FA_out_2652}=REGS_1326+REGS_1425+REGS_1446;
  assign {FA_cout_2653,FA_out_2653}=REGS_1329+REGS_1348+REGS_1471;
  assign {FA_cout_2654,FA_out_2654}=REGS_1332+REGS_1453+REGS_1474;
  assign {FA_cout_2655,FA_out_2655}=REGS_1335+REGS_1354+REGS_1455;
  assign {FA_cout_2656,FA_out_2656}=REGS_1337+REGS_1378+REGS_1497;
  assign {FA_cout_2657,FA_out_2657}=REGS_1340+REGS_1463+REGS_1500;
  assign {FA_cout_2658,FA_out_2658}=REGS_1343+REGS_1384+REGS_1465;
  assign {FA_cout_2659,FA_out_2659}=REGS_1346+REGS_1447+REGS_1468;
  assign {FA_cout_2660,FA_out_2660}=REGS_1349+REGS_1390+REGS_1509;
  assign {FA_cout_2661,FA_out_2661}=REGS_1352+REGS_1475+REGS_1512;
  assign {FA_cout_2662,FA_out_2662}=REGS_1355+REGS_1396+REGS_1477;
  assign {FA_cout_2663,FA_out_2663}=REGS_1379+REGS_1416+REGS_1534;
  assign {FA_cout_2664,FA_out_2664}=REGS_1382+REGS_1501+REGS_1537;
  assign {FA_cout_2665,FA_out_2665}=REGS_1385+REGS_1422+REGS_1503;
  assign {FA_cout_2666,FA_out_2666}=REGS_1388+REGS_1469+REGS_1506;
  assign {FA_cout_2667,FA_out_2667}=REGS_1391+REGS_1428+REGS_1546;
  assign {FA_cout_2668,FA_out_2668}=REGS_1394+REGS_1513+REGS_1549;
  assign {FA_cout_2669,FA_out_2669}=REGS_1397+REGS_1434+REGS_1515;
  assign {FA_cout_2670,FA_out_2670}=REGS_1402+REGS_1482+REGS_1518;
  assign {FA_cout_2671,FA_out_2671}=REGS_1403+REGS_1483+REGS_1519;
  assign {FA_cout_2672,FA_out_2672}=REGS_1404+REGS_1484+REGS_1520;
  assign {FA_cout_2673,FA_out_2673}=REGS_1405+REGS_1485+REGS_1521;
  assign {FA_cout_2674,FA_out_2674}=REGS_1406+REGS_1486+REGS_1522;
  assign {FA_cout_2675,FA_out_2675}=REGS_1407+REGS_1487+REGS_1523;
  assign {FA_cout_2676,FA_out_2676}=REGS_1408+REGS_1488+REGS_1524;
  assign {FA_cout_2677,FA_out_2677}=REGS_1409+REGS_1489+REGS_1525;
  assign {FA_cout_2678,FA_out_2678}=REGS_1410+REGS_1490+REGS_1526;
  assign {FA_cout_2679,FA_out_2679}=REGS_1411+REGS_1491+REGS_1527;
  assign {FA_cout_2680,FA_out_2680}=REGS_1412+REGS_1492+REGS_1528;
  assign {FA_cout_2681,FA_out_2681}=REGS_1413+REGS_1493+REGS_1529;
  assign {FA_cout_2682,FA_out_2682}=REGS_1414+REGS_1494+REGS_1530;
  assign {FA_cout_2683,FA_out_2683}=REGS_1415+REGS_1495+REGS_1531;
  assign {FA_cout_2684,FA_out_2684}=REGS_1417+REGS_1438+REGS_1558;
  assign {FA_cout_2685,FA_out_2685}=REGS_1420+REGS_1538+REGS_1561;
  assign {FA_cout_2686,FA_out_2686}=REGS_1423+REGS_1444+REGS_1540;
  assign {FA_cout_2687,FA_out_2687}=REGS_1426+REGS_1507+REGS_1543;
  assign {FA_cout_2688,FA_out_2688}=REGS_1429+REGS_1450+REGS_1570;
  assign {FA_cout_2689,FA_out_2689}=REGS_1432+REGS_1550+REGS_1573;
  assign {FA_cout_2690,FA_out_2690}=REGS_1435+REGS_1456+REGS_1552;
  assign {FA_cout_2691,FA_out_2691}=REGS_1436+REGS_1532+REGS_1555;
  assign {FA_cout_2692,FA_out_2692}=REGS_1439+REGS_1460+REGS_1582;
  assign {FA_cout_2693,FA_out_2693}=REGS_1442+REGS_1562+REGS_1585;
  assign {FA_cout_2694,FA_out_2694}=REGS_1445+REGS_1466+REGS_1564;
  assign {FA_cout_2695,FA_out_2695}=REGS_1448+REGS_1544+REGS_1567;
  assign {FA_cout_2696,FA_out_2696}=REGS_1451+REGS_1472+REGS_1594;
  assign {FA_cout_2697,FA_out_2697}=REGS_1454+REGS_1574+REGS_1597;
  assign {FA_cout_2698,FA_out_2698}=REGS_1457+REGS_1478+REGS_1576;
  assign {FA_cout_2699,FA_out_2699}=REGS_1458+REGS_1556+REGS_1579;
  assign {FA_cout_2700,FA_out_2700}=REGS_1461+REGS_1498+REGS_1606;
  assign {FA_cout_2701,FA_out_2701}=REGS_1464+REGS_1586+REGS_1609;
  assign {FA_cout_2702,FA_out_2702}=REGS_1467+REGS_1504+REGS_1588;
  assign {FA_cout_2703,FA_out_2703}=REGS_1470+REGS_1568+REGS_1591;
  assign {FA_cout_2704,FA_out_2704}=REGS_1473+REGS_1510+REGS_1618;
  assign {FA_cout_2705,FA_out_2705}=REGS_1476+REGS_1598+REGS_1621;
  assign {FA_cout_2706,FA_out_2706}=REGS_1479+REGS_1516+REGS_1600;
  assign {FA_cout_2707,FA_out_2707}=REGS_1496+REGS_1580+REGS_1603;
  assign {FA_cout_2708,FA_out_2708}=REGS_1499+REGS_1535+REGS_1643;
  assign {FA_cout_2709,FA_out_2709}=REGS_1502+REGS_1610+REGS_1646;
  assign {FA_cout_2710,FA_out_2710}=REGS_1505+REGS_1541+REGS_1612;
  assign {FA_cout_2711,FA_out_2711}=REGS_1508+REGS_1592+REGS_1615;
  assign {FA_cout_2712,FA_out_2712}=REGS_1511+REGS_1547+REGS_1655;
  assign {FA_cout_2713,FA_out_2713}=REGS_1514+REGS_1622+REGS_1658;
  assign {FA_cout_2714,FA_out_2714}=REGS_1517+REGS_1553+REGS_1624;
  assign {FA_cout_2715,FA_out_2715}=REGS_1533+REGS_1604+REGS_1640;
  assign {FA_cout_2716,FA_out_2716}=REGS_1536+REGS_1559+REGS_1676;
  assign {FA_cout_2717,FA_out_2717}=REGS_1539+REGS_1647+REGS_1679;
  assign {FA_cout_2718,FA_out_2718}=REGS_1542+REGS_1565+REGS_1649;
  assign {FA_cout_2719,FA_out_2719}=REGS_1545+REGS_1616+REGS_1652;
  assign {FA_cout_2720,FA_out_2720}=REGS_1548+REGS_1571+REGS_1688;
  assign {FA_cout_2721,FA_out_2721}=REGS_1551+REGS_1659+REGS_1691;
  assign {FA_cout_2722,FA_out_2722}=REGS_1554+REGS_1577+REGS_1661;
  assign {FA_cout_2723,FA_out_2723}=REGS_1557+REGS_1641+REGS_1673;
  assign {FA_cout_2724,FA_out_2724}=REGS_1560+REGS_1583+REGS_1702;
  assign {FA_cout_2725,FA_out_2725}=REGS_1563+REGS_1680+REGS_1705;
  assign {FA_cout_2726,FA_out_2726}=REGS_1566+REGS_1589+REGS_1682;
  assign {FA_cout_2727,FA_out_2727}=REGS_1569+REGS_1653+REGS_1685;
  assign {FA_cout_2728,FA_out_2728}=REGS_1572+REGS_1595+REGS_1714;
  assign {FA_cout_2729,FA_out_2729}=REGS_1575+REGS_1692+REGS_1717;
  assign {FA_cout_2730,FA_out_2730}=REGS_1578+REGS_1601+REGS_1694;
  assign {FA_cout_2731,FA_out_2731}=REGS_1581+REGS_1674+REGS_1699;
  assign {FA_cout_2732,FA_out_2732}=REGS_1584+REGS_1607+REGS_1728;
  assign {FA_cout_2733,FA_out_2733}=REGS_1587+REGS_1706+REGS_1731;
  assign {FA_cout_2734,FA_out_2734}=REGS_1590+REGS_1613+REGS_1708;
  assign {FA_cout_2735,FA_out_2735}=REGS_1593+REGS_1686+REGS_1711;
  assign {FA_cout_2736,FA_out_2736}=REGS_1596+REGS_1619+REGS_1740;
  assign {FA_cout_2737,FA_out_2737}=REGS_1599+REGS_1718+REGS_1743;
  assign {FA_cout_2738,FA_out_2738}=REGS_1602+REGS_1625+REGS_1720;
  assign {FA_cout_2739,FA_out_2739}=REGS_1605+REGS_1700+REGS_1725;
  assign {FA_cout_2740,FA_out_2740}=REGS_1608+REGS_1644+REGS_1761;
  assign {FA_cout_2741,FA_out_2741}=REGS_1611+REGS_1732+REGS_1764;
  assign {FA_cout_2742,FA_out_2742}=REGS_1614+REGS_1650+REGS_1734;
  assign {FA_cout_2743,FA_out_2743}=REGS_1617+REGS_1712+REGS_1737;
  assign {FA_cout_2744,FA_out_2744}=REGS_1620+REGS_1656+REGS_1773;
  assign {FA_cout_2745,FA_out_2745}=REGS_1623+REGS_1744+REGS_1776;
  assign {FA_cout_2746,FA_out_2746}=REGS_1626+REGS_1662+REGS_1746;
  assign {FA_cout_2747,FA_out_2747}=REGS_1632+REGS_1666+REGS_1749;
  assign {FA_cout_2748,FA_out_2748}=REGS_1633+REGS_1667+REGS_1750;
  assign {FA_cout_2749,FA_out_2749}=REGS_1634+REGS_1668+REGS_1751;
  assign {FA_cout_2750,FA_out_2750}=REGS_1635+REGS_1669+REGS_1752;
  assign {FA_cout_2751,FA_out_2751}=REGS_1636+REGS_1670+REGS_1753;
  assign {FA_cout_2752,FA_out_2752}=REGS_1637+REGS_1671+REGS_1754;
  assign {FA_cout_2753,FA_out_2753}=REGS_1638+REGS_1672+REGS_1755;
  assign {FA_cout_2754,FA_out_2754}=REGS_1639+REGS_1697+REGS_1787;
  assign {FA_cout_2755,FA_out_2755}=REGS_1642+REGS_1726+REGS_1758;
  assign {FA_cout_2756,FA_out_2756}=REGS_1645+REGS_1677+REGS_1793;
  assign {FA_cout_2757,FA_out_2757}=REGS_1648+REGS_1765+REGS_1796;
  assign {FA_cout_2758,FA_out_2758}=REGS_1651+REGS_1683+REGS_1767;
  assign {FA_cout_2759,FA_out_2759}=REGS_1654+REGS_1738+REGS_1770;
  assign {FA_cout_2760,FA_out_2760}=REGS_1657+REGS_1689+REGS_1805;
  assign {FA_cout_2761,FA_out_2761}=REGS_1660+REGS_1777+REGS_1808;
  assign {FA_cout_2762,FA_out_2762}=REGS_1663+REGS_1695+REGS_1779;
  assign {FA_cout_2763,FA_out_2763}=REGS_1675+REGS_1759+REGS_1790;
  assign {FA_cout_2764,FA_out_2764}=REGS_1678+REGS_1703+REGS_1821;
  assign {FA_cout_2765,FA_out_2765}=REGS_1681+REGS_1797+REGS_1824;
  assign {FA_cout_2766,FA_out_2766}=REGS_1684+REGS_1709+REGS_1799;
  assign {FA_cout_2767,FA_out_2767}=REGS_1687+REGS_1771+REGS_1802;
  assign {FA_cout_2768,FA_out_2768}=REGS_1690+REGS_1715+REGS_1833;
  assign {FA_cout_2769,FA_out_2769}=REGS_1693+REGS_1809+REGS_1836;
  assign {FA_cout_2770,FA_out_2770}=REGS_1696+REGS_1721+REGS_1811;
  assign {FA_cout_2771,FA_out_2771}=REGS_1698+REGS_1723+REGS_1815;
  assign {FA_cout_2772,FA_out_2772}=REGS_1701+REGS_1791+REGS_1818;
  assign {FA_cout_2773,FA_out_2773}=REGS_1704+REGS_1729+REGS_1847;
  assign {FA_cout_2774,FA_out_2774}=REGS_1707+REGS_1825+REGS_1849;
  assign {FA_cout_2775,FA_out_2775}=REGS_1710+REGS_1735+REGS_1827;
  assign {FA_cout_2776,FA_out_2776}=REGS_1713+REGS_1803+REGS_1830;
  assign {FA_cout_2777,FA_out_2777}=REGS_1716+REGS_1741+REGS_1856;
  assign {FA_cout_2778,FA_out_2778}=REGS_1719+REGS_1837+REGS_1858;
  assign {FA_cout_2779,FA_out_2779}=REGS_1722+REGS_1747+REGS_1839;
  assign {FA_cout_2780,FA_out_2780}=REGS_1724+REGS_1756+REGS_1863;
  assign {FA_cout_2781,FA_out_2781}=REGS_1727+REGS_1819+REGS_1845;
  assign {FA_cout_2782,FA_out_2782}=REGS_1730+REGS_1762+REGS_1868;
  assign {FA_cout_2783,FA_out_2783}=REGS_1733+REGS_1850+REGS_1870;
  assign {FA_cout_2784,FA_out_2784}=REGS_1736+REGS_1768+REGS_1872;
  assign {FA_cout_2785,FA_out_2785}=REGS_1739+REGS_1831+REGS_1854;
  assign {FA_cout_2786,FA_out_2786}=REGS_1742+REGS_1774+REGS_1877;
  assign {FA_cout_2787,FA_out_2787}=REGS_1745+REGS_1859+REGS_1879;
  assign {FA_cout_2788,FA_out_2788}=REGS_1748+REGS_1780+REGS_1881;
  assign {FA_cout_2789,FA_out_2789}=REGS_1757+REGS_1788+REGS_1886;
  assign {FA_cout_2790,FA_out_2790}=REGS_1769+REGS_1800+REGS_1889;
  assign {FA_cout_2791,FA_out_2791}=REGS_1781+REGS_1812+REGS_1892;
  assign {FA_cout_2792,FA_out_2792}=FA_cout_2206+FA_out_2207+REGS_197;
  assign {FA_cout_2793,FA_out_2793}=FA_cout_2207+FA_out_2208+REGS_198;
  assign {FA_cout_2794,FA_out_2794}=FA_cout_2208+FA_out_2209+HA_out_87;
  assign {FA_cout_2795,FA_out_2795}=FA_cout_2209+FA_out_2210+HA_cout_87;
  assign {FA_cout_2796,FA_out_2796}=FA_cout_2210+FA_out_2211+HA_cout_88;
  assign {FA_cout_2797,FA_out_2797}=FA_cout_2211+FA_out_2212+HA_cout_89;
  assign {FA_cout_2798,FA_out_2798}=FA_cout_2212+FA_out_2213+FA_cout_2270;
  assign {FA_cout_2799,FA_out_2799}=FA_cout_2213+FA_out_2214+FA_cout_2271;
  assign {FA_cout_2800,FA_out_2800}=FA_cout_2214+FA_out_2215+FA_cout_2272;
  assign {FA_cout_2801,FA_out_2801}=FA_cout_2215+FA_out_2216+FA_cout_2273;
  assign {FA_cout_2802,FA_out_2802}=FA_cout_2216+FA_out_2217+FA_cout_2274;
  assign {FA_cout_2803,FA_out_2803}=FA_cout_2217+FA_out_2218+FA_cout_2275;
  assign {FA_cout_2804,FA_out_2804}=FA_cout_2218+FA_out_2219+FA_cout_2276;
  assign {FA_cout_2805,FA_out_2805}=FA_cout_2219+FA_out_2220+FA_cout_2277;
  assign {FA_cout_2806,FA_out_2806}=FA_cout_2220+FA_out_2221+FA_cout_2278;
  assign {FA_cout_2807,FA_out_2807}=FA_cout_2221+FA_out_2222+FA_cout_2279;
  assign {FA_cout_2808,FA_out_2808}=FA_cout_2222+FA_out_2223+FA_cout_2280;
  assign {FA_cout_2809,FA_out_2809}=FA_cout_2223+FA_out_2224+FA_cout_2281;
  assign {FA_cout_2810,FA_out_2810}=FA_cout_2224+FA_out_2225+FA_cout_2282;
  assign {FA_cout_2811,FA_out_2811}=FA_cout_2225+FA_out_2226+FA_cout_2283;
  assign {FA_cout_2812,FA_out_2812}=FA_cout_2226+FA_out_2227+FA_cout_2284;
  assign {FA_cout_2813,FA_out_2813}=FA_cout_2227+FA_out_2228+FA_cout_2285;
  assign {FA_cout_2814,FA_out_2814}=FA_cout_2228+FA_out_2229+FA_cout_2286;
  assign {FA_cout_2815,FA_out_2815}=FA_cout_2229+FA_out_2230+FA_cout_2287;
  assign {FA_cout_2816,FA_out_2816}=FA_cout_2230+FA_out_2231+FA_cout_2288;
  assign {FA_cout_2817,FA_out_2817}=FA_cout_2231+FA_out_2232+FA_cout_2289;
  assign {FA_cout_2818,FA_out_2818}=FA_cout_2232+FA_out_2233+FA_cout_2290;
  assign {FA_cout_2819,FA_out_2819}=FA_cout_2233+FA_out_2234+FA_cout_2291;
  assign {FA_cout_2820,FA_out_2820}=FA_cout_2234+FA_out_2235+FA_cout_2292;
  assign {FA_cout_2821,FA_out_2821}=FA_cout_2235+FA_out_2236+FA_cout_2293;
  assign {FA_cout_2822,FA_out_2822}=FA_cout_2236+FA_out_2237+FA_cout_2294;
  assign {FA_cout_2823,FA_out_2823}=FA_cout_2237+FA_out_2238+FA_cout_2295;
  assign {FA_cout_2824,FA_out_2824}=FA_cout_2238+FA_out_2239+FA_cout_2296;
  assign {FA_cout_2825,FA_out_2825}=FA_cout_2239+FA_out_2240+FA_cout_2297;
  assign {FA_cout_2826,FA_out_2826}=FA_cout_2240+FA_out_2241+FA_cout_2298;
  assign {FA_cout_2827,FA_out_2827}=FA_cout_2241+FA_out_2242+FA_cout_2299;
  assign {FA_cout_2828,FA_out_2828}=FA_cout_2242+FA_out_2243+FA_cout_2300;
  assign {FA_cout_2829,FA_out_2829}=FA_cout_2243+FA_out_2244+FA_cout_2301;
  assign {FA_cout_2830,FA_out_2830}=FA_cout_2244+FA_out_2245+FA_cout_2302;
  assign {FA_cout_2831,FA_out_2831}=FA_cout_2245+FA_out_2246+FA_cout_2303;
  assign {FA_cout_2832,FA_out_2832}=FA_cout_2246+FA_out_2247+FA_cout_2304;
  assign {FA_cout_2833,FA_out_2833}=FA_cout_2247+FA_out_2248+FA_cout_2305;
  assign {FA_cout_2834,FA_out_2834}=FA_cout_2248+FA_out_2249+FA_cout_2306;
  assign {FA_cout_2835,FA_out_2835}=FA_cout_2249+FA_out_2250+FA_cout_2307;
  assign {FA_cout_2836,FA_out_2836}=FA_cout_2250+FA_out_2251+FA_cout_2308;
  assign {FA_cout_2837,FA_out_2837}=FA_cout_2251+FA_out_2252+FA_cout_2309;
  assign {FA_cout_2838,FA_out_2838}=FA_cout_2252+FA_out_2253+FA_cout_2310;
  assign {FA_cout_2839,FA_out_2839}=FA_cout_2253+FA_out_2254+FA_cout_2311;
  assign {FA_cout_2840,FA_out_2840}=FA_cout_2254+FA_out_2255+FA_cout_2312;
  assign {FA_cout_2841,FA_out_2841}=FA_cout_2255+FA_out_2256+FA_cout_2313;
  assign {FA_cout_2842,FA_out_2842}=FA_cout_2256+FA_out_2257+FA_cout_2314;
  assign {FA_cout_2843,FA_out_2843}=FA_cout_2257+FA_out_2258+FA_cout_2315;
  assign {FA_cout_2844,FA_out_2844}=FA_cout_2258+FA_out_2259+FA_cout_2316;
  assign {FA_cout_2845,FA_out_2845}=FA_cout_2259+FA_out_2260+FA_cout_2317;
  assign {FA_cout_2846,FA_out_2846}=FA_cout_2260+FA_out_2261+FA_cout_2318;
  assign {FA_cout_2847,FA_out_2847}=FA_cout_2261+FA_out_2262+FA_cout_2319;
  assign {FA_cout_2848,FA_out_2848}=FA_cout_2262+FA_out_2263+FA_cout_2320;
  assign {FA_cout_2849,FA_out_2849}=FA_cout_2263+FA_out_2264+FA_cout_2321;
  assign {FA_cout_2850,FA_out_2850}=FA_cout_2264+FA_out_2265+FA_cout_2322;
  assign {FA_cout_2851,FA_out_2851}=FA_cout_2265+FA_out_2266+FA_cout_2323;
  assign {FA_cout_2852,FA_out_2852}=FA_cout_2266+FA_out_2267+FA_cout_2325;
  assign {FA_cout_2853,FA_out_2853}=FA_cout_2267+FA_out_2268+FA_cout_2327;
  assign {FA_cout_2854,FA_out_2854}=FA_cout_2268+FA_out_2269+FA_cout_2329;
  assign {FA_cout_2855,FA_out_2855}=FA_cout_2269+FA_out_2324+FA_cout_2331;
  assign {FA_cout_2856,FA_out_2856}=FA_cout_2324+FA_out_2326+FA_cout_2333;
  assign {FA_cout_2857,FA_out_2857}=FA_out_2275+HA_cout_90+HA_out_91;
  assign {FA_cout_2858,FA_out_2858}=FA_out_2276+HA_cout_91+FA_out_2339;
  assign {FA_cout_2859,FA_out_2859}=FA_out_2277+FA_cout_2339+FA_out_2340;
  assign {FA_cout_2860,FA_out_2860}=FA_out_2278+FA_cout_2340+FA_out_2341;
  assign {FA_cout_2861,FA_out_2861}=FA_out_2279+FA_cout_2341+FA_out_2342;
  assign {FA_cout_2862,FA_out_2862}=FA_out_2280+FA_cout_2342+FA_out_2343;
  assign {FA_cout_2863,FA_out_2863}=FA_out_2281+FA_cout_2343+FA_out_2344;
  assign {FA_cout_2864,FA_out_2864}=FA_out_2282+FA_cout_2344+FA_out_2345;
  assign {FA_cout_2865,FA_out_2865}=FA_out_2283+FA_cout_2345+FA_out_2346;
  assign {FA_cout_2866,FA_out_2866}=FA_out_2284+FA_cout_2346+FA_out_2347;
  assign {FA_cout_2867,FA_out_2867}=FA_out_2285+FA_cout_2347+FA_out_2348;
  assign {FA_cout_2868,FA_out_2868}=FA_out_2286+FA_cout_2348+FA_out_2349;
  assign {FA_cout_2869,FA_out_2869}=FA_out_2287+FA_cout_2349+FA_out_2350;
  assign {FA_cout_2870,FA_out_2870}=FA_out_2288+FA_cout_2350+FA_out_2351;
  assign {FA_cout_2871,FA_out_2871}=FA_out_2289+FA_cout_2351+FA_out_2352;
  assign {FA_cout_2872,FA_out_2872}=FA_out_2290+FA_cout_2352+FA_out_2353;
  assign {FA_cout_2873,FA_out_2873}=FA_out_2291+FA_cout_2353+FA_out_2354;
  assign {FA_cout_2874,FA_out_2874}=FA_out_2292+FA_cout_2354+FA_out_2355;
  assign {FA_cout_2875,FA_out_2875}=FA_out_2293+FA_cout_2355+FA_out_2356;
  assign {FA_cout_2876,FA_out_2876}=FA_out_2294+FA_cout_2356+FA_out_2357;
  assign {FA_cout_2877,FA_out_2877}=FA_out_2295+FA_cout_2357+FA_out_2358;
  assign {FA_cout_2878,FA_out_2878}=FA_out_2296+FA_cout_2358+FA_out_2359;
  assign {FA_cout_2879,FA_out_2879}=FA_out_2297+FA_cout_2359+FA_out_2360;
  assign {FA_cout_2880,FA_out_2880}=FA_out_2298+FA_cout_2360+FA_out_2361;
  assign {FA_cout_2881,FA_out_2881}=FA_out_2299+FA_cout_2361+FA_out_2362;
  assign {FA_cout_2882,FA_out_2882}=FA_out_2300+FA_cout_2362+FA_out_2363;
  assign {FA_cout_2883,FA_out_2883}=FA_out_2301+FA_cout_2363+FA_out_2364;
  assign {FA_cout_2884,FA_out_2884}=FA_out_2302+FA_cout_2364+FA_out_2365;
  assign {FA_cout_2885,FA_out_2885}=FA_out_2303+FA_cout_2365+FA_out_2366;
  assign {FA_cout_2886,FA_out_2886}=FA_out_2304+FA_cout_2366+FA_out_2367;
  assign {FA_cout_2887,FA_out_2887}=FA_out_2305+FA_cout_2367+FA_out_2368;
  assign {FA_cout_2888,FA_out_2888}=FA_out_2306+FA_cout_2368+FA_out_2369;
  assign {FA_cout_2889,FA_out_2889}=FA_out_2307+FA_cout_2369+FA_out_2370;
  assign {FA_cout_2890,FA_out_2890}=FA_out_2308+FA_cout_2370+FA_out_2371;
  assign {FA_cout_2891,FA_out_2891}=FA_out_2309+FA_cout_2371+FA_out_2372;
  assign {FA_cout_2892,FA_out_2892}=FA_out_2310+FA_cout_2372+FA_out_2373;
  assign {FA_cout_2893,FA_out_2893}=FA_out_2311+FA_cout_2373+FA_out_2374;
  assign {FA_cout_2894,FA_out_2894}=FA_out_2312+FA_cout_2374+FA_out_2375;
  assign {FA_cout_2895,FA_out_2895}=FA_out_2313+FA_cout_2375+FA_out_2376;
  assign {FA_cout_2896,FA_out_2896}=FA_out_2314+FA_cout_2376+FA_out_2377;
  assign {FA_cout_2897,FA_out_2897}=FA_out_2315+FA_cout_2377+FA_out_2378;
  assign {FA_cout_2898,FA_out_2898}=FA_out_2316+FA_cout_2378+FA_out_2379;
  assign {FA_cout_2899,FA_out_2899}=FA_out_2317+FA_cout_2379+FA_out_2380;
  assign {FA_cout_2900,FA_out_2900}=FA_out_2318+FA_cout_2380+FA_out_2381;
  assign {FA_cout_2901,FA_out_2901}=FA_out_2319+FA_cout_2381+FA_out_2382;
  assign {FA_cout_2902,FA_out_2902}=FA_out_2320+FA_cout_2382+FA_out_2383;
  assign {FA_cout_2903,FA_out_2903}=FA_out_2321+FA_cout_2383+FA_out_2384;
  assign {FA_cout_2904,FA_out_2904}=FA_out_2322+FA_cout_2384+FA_out_2385;
  assign {FA_cout_2905,FA_out_2905}=FA_out_2323+FA_cout_2385+FA_out_2386;
  assign {FA_cout_2906,FA_out_2906}=FA_out_2325+FA_cout_2386+FA_out_2389;
  assign {FA_cout_2907,FA_out_2907}=FA_cout_2326+FA_out_2328+FA_cout_2335;
  assign {FA_cout_2908,FA_out_2908}=FA_out_2327+FA_cout_2389+FA_out_2392;
  assign {FA_cout_2909,FA_out_2909}=FA_cout_2328+FA_out_2330+FA_cout_2337;
  assign {FA_cout_2910,FA_out_2910}=FA_out_2329+FA_cout_2392+FA_out_2395;
  assign {FA_cout_2911,FA_out_2911}=FA_cout_2330+FA_out_2332+FA_cout_2387;
  assign {FA_cout_2912,FA_out_2912}=FA_out_2331+FA_cout_2395+FA_out_2398;
  assign {FA_cout_2913,FA_out_2913}=FA_cout_2332+FA_out_2334+FA_cout_2390;
  assign {FA_cout_2914,FA_out_2914}=FA_out_2333+FA_cout_2398+FA_out_2401;
  assign {FA_cout_2915,FA_out_2915}=FA_cout_2334+FA_out_2336+FA_cout_2393;
  assign {FA_cout_2916,FA_out_2916}=FA_out_2335+FA_cout_2401+FA_out_2445;
  assign {FA_cout_2917,FA_out_2917}=FA_cout_2336+FA_out_2338+FA_cout_2396;
  assign {FA_cout_2918,FA_out_2918}=FA_out_2337+FA_cout_2445+FA_out_2449;
  assign {FA_cout_2919,FA_out_2919}=FA_cout_2338+FA_out_2388+FA_cout_2399;
  assign {FA_cout_2920,FA_out_2920}=FA_out_2387+FA_cout_2449+FA_out_2453;
  assign {FA_cout_2921,FA_out_2921}=FA_cout_2388+FA_out_2391+FA_cout_2402;
  assign {FA_cout_2922,FA_out_2922}=FA_out_2390+FA_cout_2453+FA_out_2457;
  assign {FA_cout_2923,FA_out_2923}=FA_cout_2391+FA_out_2394+FA_cout_2446;
  assign {FA_cout_2924,FA_out_2924}=FA_out_2393+FA_cout_2457+FA_out_2461;
  assign {FA_cout_2925,FA_out_2925}=FA_cout_2394+FA_out_2397+FA_cout_2450;
  assign {FA_cout_2926,FA_out_2926}=FA_out_2396+FA_cout_2461+FA_out_2465;
  assign {FA_cout_2927,FA_out_2927}=FA_cout_2397+FA_out_2400+FA_cout_2454;
  assign {FA_cout_2928,FA_out_2928}=FA_out_2399+FA_cout_2465+FA_out_2469;
  assign {FA_cout_2929,FA_out_2929}=FA_cout_2400+FA_out_2403+FA_cout_2458;
  assign {FA_cout_2930,FA_out_2930}=FA_out_2402+FA_cout_2469+FA_out_2473;
  assign {FA_cout_2931,FA_out_2931}=FA_cout_2403+FA_out_2447+FA_cout_2462;
  assign {FA_cout_2932,FA_out_2932}=FA_cout_2405+FA_out_2406+REGS_813;
  assign {FA_cout_2933,FA_out_2933}=FA_cout_2406+FA_out_2407+REGS_814;
  assign {FA_cout_2934,FA_out_2934}=FA_cout_2407+FA_out_2408+REGS_815;
  assign {FA_cout_2935,FA_out_2935}=FA_cout_2408+FA_out_2409+HA_out_94;
  assign {FA_cout_2936,FA_out_2936}=FA_cout_2409+FA_out_2410+HA_cout_94;
  assign {FA_cout_2937,FA_out_2937}=FA_cout_2410+FA_out_2411+HA_cout_95;
  assign {FA_cout_2938,FA_out_2938}=FA_cout_2411+FA_out_2412+FA_cout_2476;
  assign {FA_cout_2939,FA_out_2939}=FA_cout_2412+FA_out_2413+FA_cout_2477;
  assign {FA_cout_2940,FA_out_2940}=FA_cout_2413+FA_out_2414+FA_cout_2478;
  assign {FA_cout_2941,FA_out_2941}=FA_cout_2414+FA_out_2415+FA_cout_2479;
  assign {FA_cout_2942,FA_out_2942}=FA_cout_2415+FA_out_2416+FA_cout_2480;
  assign {FA_cout_2943,FA_out_2943}=FA_cout_2416+FA_out_2417+FA_cout_2481;
  assign {FA_cout_2944,FA_out_2944}=FA_cout_2417+FA_out_2418+FA_cout_2482;
  assign {FA_cout_2945,FA_out_2945}=FA_cout_2418+FA_out_2419+FA_cout_2483;
  assign {FA_cout_2946,FA_out_2946}=FA_cout_2419+FA_out_2420+FA_cout_2484;
  assign {FA_cout_2947,FA_out_2947}=FA_cout_2420+FA_out_2421+FA_cout_2485;
  assign {FA_cout_2948,FA_out_2948}=FA_cout_2421+FA_out_2422+FA_cout_2486;
  assign {FA_cout_2949,FA_out_2949}=FA_cout_2422+FA_out_2423+FA_cout_2487;
  assign {FA_cout_2950,FA_out_2950}=FA_cout_2423+FA_out_2424+FA_cout_2488;
  assign {FA_cout_2951,FA_out_2951}=FA_cout_2424+FA_out_2425+FA_cout_2489;
  assign {FA_cout_2952,FA_out_2952}=FA_cout_2425+FA_out_2426+FA_cout_2490;
  assign {FA_cout_2953,FA_out_2953}=FA_cout_2426+FA_out_2427+FA_cout_2491;
  assign {FA_cout_2954,FA_out_2954}=FA_cout_2427+FA_out_2428+FA_cout_2492;
  assign {FA_cout_2955,FA_out_2955}=FA_cout_2428+FA_out_2429+FA_cout_2493;
  assign {FA_cout_2956,FA_out_2956}=FA_cout_2429+FA_out_2430+FA_cout_2494;
  assign {FA_cout_2957,FA_out_2957}=FA_cout_2430+FA_out_2431+FA_cout_2495;
  assign {FA_cout_2958,FA_out_2958}=FA_cout_2431+FA_out_2432+FA_cout_2496;
  assign {FA_cout_2959,FA_out_2959}=FA_cout_2432+FA_out_2433+FA_cout_2497;
  assign {FA_cout_2960,FA_out_2960}=FA_cout_2433+FA_out_2434+FA_cout_2498;
  assign {FA_cout_2961,FA_out_2961}=FA_cout_2434+FA_out_2435+FA_cout_2499;
  assign {FA_cout_2962,FA_out_2962}=FA_cout_2435+FA_out_2436+FA_cout_2500;
  assign {FA_cout_2963,FA_out_2963}=FA_cout_2436+FA_out_2437+FA_cout_2501;
  assign {FA_cout_2964,FA_out_2964}=FA_cout_2437+FA_out_2438+FA_cout_2502;
  assign {FA_cout_2965,FA_out_2965}=FA_cout_2438+FA_out_2439+FA_cout_2503;
  assign {FA_cout_2966,FA_out_2966}=FA_cout_2439+FA_out_2440+FA_cout_2504;
  assign {FA_cout_2967,FA_out_2967}=FA_cout_2440+FA_out_2441+FA_cout_2505;
  assign {FA_cout_2968,FA_out_2968}=FA_cout_2441+FA_out_2442+FA_cout_2506;
  assign {FA_cout_2969,FA_out_2969}=FA_cout_2442+FA_out_2443+FA_cout_2507;
  assign {FA_cout_2970,FA_out_2970}=FA_cout_2443+FA_out_2444+FA_cout_2508;
  assign {FA_cout_2971,FA_out_2971}=FA_cout_2444+FA_out_2448+FA_cout_2509;
  assign {FA_cout_2972,FA_out_2972}=FA_out_2446+FA_cout_2473+FA_out_2512;
  assign {FA_cout_2973,FA_out_2973}=FA_cout_2447+FA_out_2451+FA_cout_2466;
  assign {FA_cout_2974,FA_out_2974}=FA_cout_2448+FA_out_2452+FA_cout_2510;
  assign {FA_cout_2975,FA_out_2975}=FA_out_2450+FA_cout_2512+FA_out_2516;
  assign {FA_cout_2976,FA_out_2976}=FA_cout_2451+FA_out_2455+FA_cout_2470;
  assign {FA_cout_2977,FA_out_2977}=FA_cout_2452+FA_out_2456+FA_cout_2519;
  assign {FA_cout_2978,FA_out_2978}=FA_out_2454+FA_cout_2516+FA_out_2521;
  assign {FA_cout_2979,FA_out_2979}=FA_cout_2455+FA_out_2459+FA_cout_2474;
  assign {FA_cout_2980,FA_out_2980}=FA_cout_2456+FA_out_2460+FA_cout_2524;
  assign {FA_cout_2981,FA_out_2981}=FA_out_2458+FA_cout_2521+FA_out_2526;
  assign {FA_cout_2982,FA_out_2982}=FA_cout_2459+FA_out_2463+FA_cout_2513;
  assign {FA_cout_2983,FA_out_2983}=FA_cout_2460+FA_out_2464+FA_cout_2529;
  assign {FA_cout_2984,FA_out_2984}=FA_out_2462+FA_cout_2526+FA_out_2531;
  assign {FA_cout_2985,FA_out_2985}=FA_cout_2463+FA_out_2467+FA_cout_2517;
  assign {FA_cout_2986,FA_out_2986}=FA_cout_2464+FA_out_2468+FA_cout_2561;
  assign {FA_cout_2987,FA_out_2987}=FA_out_2466+FA_cout_2531+FA_out_2563;
  assign {FA_cout_2988,FA_out_2988}=FA_cout_2467+FA_out_2471+FA_cout_2522;
  assign {FA_cout_2989,FA_out_2989}=FA_cout_2468+FA_out_2472+FA_cout_2567;
  assign {FA_cout_2990,FA_out_2990}=FA_out_2470+FA_cout_2563+FA_out_2569;
  assign {FA_cout_2991,FA_out_2991}=FA_cout_2471+FA_out_2475+FA_cout_2527;
  assign {FA_cout_2992,FA_out_2992}=FA_cout_2472+FA_out_2511+FA_cout_2573;
  assign {FA_cout_2993,FA_out_2993}=FA_out_2474+FA_cout_2569+FA_out_2575;
  assign {FA_cout_2994,FA_out_2994}=FA_cout_2475+FA_out_2514+FA_cout_2532;
  assign {FA_cout_2995,FA_out_2995}=FA_cout_2511+FA_out_2515+FA_cout_2579;
  assign {FA_cout_2996,FA_out_2996}=FA_out_2513+FA_cout_2575+FA_out_2581;
  assign {FA_cout_2997,FA_out_2997}=FA_cout_2514+FA_out_2518+FA_cout_2564;
  assign {FA_cout_2998,FA_out_2998}=FA_out_2481+HA_cout_96+HA_out_97;
  assign {FA_cout_2999,FA_out_2999}=FA_out_2482+HA_cout_97+HA_out_98;
  assign {FA_cout_3000,FA_out_3000}=FA_out_2483+HA_cout_98+FA_out_2534;
  assign {FA_cout_3001,FA_out_3001}=FA_out_2484+FA_cout_2534+FA_out_2535;
  assign {FA_cout_3002,FA_out_3002}=FA_out_2485+FA_cout_2535+FA_out_2536;
  assign {FA_cout_3003,FA_out_3003}=FA_out_2486+FA_cout_2536+FA_out_2537;
  assign {FA_cout_3004,FA_out_3004}=FA_out_2487+FA_cout_2537+FA_out_2538;
  assign {FA_cout_3005,FA_out_3005}=FA_out_2488+FA_cout_2538+FA_out_2539;
  assign {FA_cout_3006,FA_out_3006}=FA_out_2489+FA_cout_2539+FA_out_2540;
  assign {FA_cout_3007,FA_out_3007}=FA_out_2490+FA_cout_2540+FA_out_2541;
  assign {FA_cout_3008,FA_out_3008}=FA_out_2491+FA_cout_2541+FA_out_2542;
  assign {FA_cout_3009,FA_out_3009}=FA_out_2492+FA_cout_2542+FA_out_2543;
  assign {FA_cout_3010,FA_out_3010}=FA_out_2493+FA_cout_2543+FA_out_2544;
  assign {FA_cout_3011,FA_out_3011}=FA_out_2494+FA_cout_2544+FA_out_2545;
  assign {FA_cout_3012,FA_out_3012}=FA_out_2495+FA_cout_2545+FA_out_2546;
  assign {FA_cout_3013,FA_out_3013}=FA_out_2496+FA_cout_2546+FA_out_2547;
  assign {FA_cout_3014,FA_out_3014}=FA_out_2497+FA_cout_2547+FA_out_2548;
  assign {FA_cout_3015,FA_out_3015}=FA_out_2498+FA_cout_2548+FA_out_2549;
  assign {FA_cout_3016,FA_out_3016}=FA_out_2499+FA_cout_2549+FA_out_2550;
  assign {FA_cout_3017,FA_out_3017}=FA_out_2500+FA_cout_2550+FA_out_2551;
  assign {FA_cout_3018,FA_out_3018}=FA_out_2501+FA_cout_2551+FA_out_2552;
  assign {FA_cout_3019,FA_out_3019}=FA_out_2502+FA_cout_2552+FA_out_2553;
  assign {FA_cout_3020,FA_out_3020}=FA_out_2503+FA_cout_2553+FA_out_2554;
  assign {FA_cout_3021,FA_out_3021}=FA_out_2504+FA_cout_2554+FA_out_2555;
  assign {FA_cout_3022,FA_out_3022}=FA_out_2505+FA_cout_2555+FA_out_2556;
  assign {FA_cout_3023,FA_out_3023}=FA_out_2506+FA_cout_2556+FA_out_2557;
  assign {FA_cout_3024,FA_out_3024}=FA_out_2507+FA_cout_2557+FA_out_2558;
  assign {FA_cout_3025,FA_out_3025}=FA_out_2508+FA_cout_2558+FA_out_2559;
  assign {FA_cout_3026,FA_out_3026}=FA_out_2509+FA_cout_2559+FA_out_2560;
  assign {FA_cout_3027,FA_out_3027}=FA_out_2510+FA_cout_2560+FA_out_2566;
  assign {FA_cout_3028,FA_out_3028}=FA_cout_2515+FA_out_2520+FA_cout_2585;
  assign {FA_cout_3029,FA_out_3029}=FA_out_2517+FA_cout_2581+FA_out_2587;
  assign {FA_cout_3030,FA_out_3030}=FA_cout_2518+FA_out_2523+FA_cout_2570;
  assign {FA_cout_3031,FA_out_3031}=FA_out_2519+FA_cout_2566+FA_out_2572;
  assign {FA_cout_3032,FA_out_3032}=FA_cout_2520+FA_out_2525+FA_cout_2591;
  assign {FA_cout_3033,FA_out_3033}=FA_out_2522+FA_cout_2587+FA_out_2593;
  assign {FA_cout_3034,FA_out_3034}=FA_cout_2523+FA_out_2528+FA_cout_2576;
  assign {FA_cout_3035,FA_out_3035}=FA_out_2524+FA_cout_2572+FA_out_2578;
  assign {FA_cout_3036,FA_out_3036}=FA_cout_2525+FA_out_2530+FA_cout_2597;
  assign {FA_cout_3037,FA_out_3037}=FA_out_2527+FA_cout_2593+FA_out_2599;
  assign {FA_cout_3038,FA_out_3038}=FA_cout_2528+FA_out_2533+FA_cout_2582;
  assign {FA_cout_3039,FA_out_3039}=FA_out_2529+FA_cout_2578+FA_out_2584;
  assign {FA_cout_3040,FA_out_3040}=FA_cout_2530+FA_out_2562+FA_cout_2603;
  assign {FA_cout_3041,FA_out_3041}=FA_out_2532+FA_cout_2599+FA_out_2605;
  assign {FA_cout_3042,FA_out_3042}=FA_cout_2533+FA_out_2565+FA_cout_2588;
  assign {FA_cout_3043,FA_out_3043}=FA_out_2561+FA_cout_2584+FA_out_2590;
  assign {FA_cout_3044,FA_out_3044}=FA_cout_2562+FA_out_2568+FA_cout_2630;
  assign {FA_cout_3045,FA_out_3045}=FA_out_2564+FA_cout_2605+FA_out_2632;
  assign {FA_cout_3046,FA_out_3046}=FA_cout_2565+FA_out_2571+FA_cout_2594;
  assign {FA_cout_3047,FA_out_3047}=FA_out_2567+FA_cout_2590+FA_out_2596;
  assign {FA_cout_3048,FA_out_3048}=FA_cout_2568+FA_out_2574+FA_cout_2637;
  assign {FA_cout_3049,FA_out_3049}=FA_out_2570+FA_cout_2632+FA_out_2639;
  assign {FA_cout_3050,FA_out_3050}=FA_cout_2571+FA_out_2577+FA_cout_2600;
  assign {FA_cout_3051,FA_out_3051}=FA_out_2573+FA_cout_2596+FA_out_2602;
  assign {FA_cout_3052,FA_out_3052}=FA_cout_2574+FA_out_2580+FA_cout_2644;
  assign {FA_cout_3053,FA_out_3053}=FA_out_2576+FA_cout_2639+FA_out_2646;
  assign {FA_cout_3054,FA_out_3054}=FA_cout_2577+FA_out_2583+FA_cout_2606;
  assign {FA_cout_3055,FA_out_3055}=FA_out_2579+FA_cout_2602+FA_out_2629;
  assign {FA_cout_3056,FA_out_3056}=FA_cout_2580+FA_out_2586+FA_cout_2651;
  assign {FA_cout_3057,FA_out_3057}=FA_out_2582+FA_cout_2646+FA_out_2653;
  assign {FA_cout_3058,FA_out_3058}=FA_cout_2583+FA_out_2589+FA_cout_2633;
  assign {FA_cout_3059,FA_out_3059}=FA_out_2585+FA_cout_2629+FA_out_2636;
  assign {FA_cout_3060,FA_out_3060}=FA_cout_2586+FA_out_2592+FA_cout_2658;
  assign {FA_cout_3061,FA_out_3061}=FA_out_2588+FA_cout_2653+FA_out_2660;
  assign {FA_cout_3062,FA_out_3062}=FA_cout_2589+FA_out_2595+FA_cout_2640;
  assign {FA_cout_3063,FA_out_3063}=FA_out_2591+FA_cout_2636+FA_out_2643;
  assign {FA_cout_3064,FA_out_3064}=FA_cout_2592+FA_out_2598+FA_cout_2665;
  assign {FA_cout_3065,FA_out_3065}=FA_out_2594+FA_cout_2660+FA_out_2667;
  assign {FA_cout_3066,FA_out_3066}=FA_cout_2595+FA_out_2601+FA_cout_2647;
  assign {FA_cout_3067,FA_out_3067}=FA_out_2597+FA_cout_2643+FA_out_2650;
  assign {FA_cout_3068,FA_out_3068}=FA_cout_2598+FA_out_2604+FA_cout_2686;
  assign {FA_cout_3069,FA_out_3069}=FA_out_2600+FA_cout_2667+FA_out_2688;
  assign {FA_cout_3070,FA_out_3070}=FA_cout_2601+FA_out_2607+FA_cout_2654;
  assign {FA_cout_3071,FA_out_3071}=FA_out_2603+FA_cout_2650+FA_out_2657;
  assign {FA_cout_3072,FA_out_3072}=FA_cout_2604+FA_out_2631+FA_cout_2694;
  assign {FA_cout_3073,FA_out_3073}=FA_out_2606+FA_cout_2688+FA_out_2696;
  assign {FA_cout_3074,FA_out_3074}=FA_cout_2607+FA_out_2634+FA_cout_2661;
  assign {FA_cout_3075,FA_out_3075}=FA_cout_2610+FA_out_2611+REGS_1398;
  assign {FA_cout_3076,FA_out_3076}=FA_cout_2611+FA_out_2612+REGS_1399;
  assign {FA_cout_3077,FA_out_3077}=FA_cout_2612+FA_out_2613+HA_out_101;
  assign {FA_cout_3078,FA_out_3078}=FA_cout_2613+FA_out_2614+HA_cout_101;
  assign {FA_cout_3079,FA_out_3079}=FA_cout_2614+FA_out_2615+HA_cout_102;
  assign {FA_cout_3080,FA_out_3080}=FA_cout_2615+FA_out_2616+FA_cout_2670;
  assign {FA_cout_3081,FA_out_3081}=FA_cout_2616+FA_out_2617+FA_cout_2671;
  assign {FA_cout_3082,FA_out_3082}=FA_cout_2617+FA_out_2618+FA_cout_2672;
  assign {FA_cout_3083,FA_out_3083}=FA_cout_2618+FA_out_2619+FA_cout_2673;
  assign {FA_cout_3084,FA_out_3084}=FA_cout_2619+FA_out_2620+FA_cout_2674;
  assign {FA_cout_3085,FA_out_3085}=FA_cout_2620+FA_out_2621+FA_cout_2675;
  assign {FA_cout_3086,FA_out_3086}=FA_cout_2621+FA_out_2622+FA_cout_2676;
  assign {FA_cout_3087,FA_out_3087}=FA_cout_2622+FA_out_2623+FA_cout_2677;
  assign {FA_cout_3088,FA_out_3088}=FA_cout_2623+FA_out_2624+FA_cout_2678;
  assign {FA_cout_3089,FA_out_3089}=FA_cout_2624+FA_out_2625+FA_cout_2679;
  assign {FA_cout_3090,FA_out_3090}=FA_cout_2625+FA_out_2626+FA_cout_2680;
  assign {FA_cout_3091,FA_out_3091}=FA_cout_2626+FA_out_2627+FA_cout_2681;
  assign {FA_cout_3092,FA_out_3092}=FA_cout_2627+FA_out_2628+FA_cout_2682;
  assign {FA_cout_3093,FA_out_3093}=FA_cout_2628+FA_out_2635+FA_cout_2683;
  assign {FA_cout_3094,FA_out_3094}=FA_out_2630+FA_cout_2657+FA_out_2664;
  assign {FA_cout_3095,FA_out_3095}=FA_cout_2631+FA_out_2638+FA_cout_2702;
  assign {FA_cout_3096,FA_out_3096}=FA_out_2633+FA_cout_2696+FA_out_2704;
  assign {FA_cout_3097,FA_out_3097}=FA_cout_2634+FA_out_2641+FA_cout_2668;
  assign {FA_cout_3098,FA_out_3098}=FA_cout_2635+FA_out_2642+FA_cout_2691;
  assign {FA_cout_3099,FA_out_3099}=FA_out_2637+FA_cout_2664+FA_out_2685;
  assign {FA_cout_3100,FA_out_3100}=FA_cout_2638+FA_out_2645+FA_cout_2710;
  assign {FA_cout_3101,FA_out_3101}=FA_out_2640+FA_cout_2704+FA_out_2712;
  assign {FA_cout_3102,FA_out_3102}=FA_cout_2641+FA_out_2648+FA_cout_2689;
  assign {FA_cout_3103,FA_out_3103}=FA_cout_2642+FA_out_2649+FA_cout_2699;
  assign {FA_cout_3104,FA_out_3104}=FA_out_2644+FA_cout_2685+FA_out_2693;
  assign {FA_cout_3105,FA_out_3105}=FA_cout_2645+FA_out_2652+FA_cout_2718;
  assign {FA_cout_3106,FA_out_3106}=FA_out_2647+FA_cout_2712+FA_out_2720;
  assign {FA_cout_3107,FA_out_3107}=FA_cout_2648+FA_out_2655+FA_cout_2697;
  assign {FA_cout_3108,FA_out_3108}=FA_cout_2649+FA_out_2656+FA_cout_2707;
  assign {FA_cout_3109,FA_out_3109}=FA_out_2651+FA_cout_2693+FA_out_2701;
  assign {FA_cout_3110,FA_out_3110}=FA_cout_2652+FA_out_2659+FA_cout_2726;
  assign {FA_cout_3111,FA_out_3111}=FA_out_2654+FA_cout_2720+FA_out_2728;
  assign {FA_cout_3112,FA_out_3112}=FA_cout_2655+FA_out_2662+FA_cout_2705;
  assign {FA_cout_3113,FA_out_3113}=FA_cout_2656+FA_out_2663+FA_cout_2715;
  assign {FA_cout_3114,FA_out_3114}=FA_out_2658+FA_cout_2701+FA_out_2709;
  assign {FA_cout_3115,FA_out_3115}=FA_cout_2659+FA_out_2666+FA_cout_2734;
  assign {FA_cout_3116,FA_out_3116}=FA_out_2661+FA_cout_2728+FA_out_2736;
  assign {FA_cout_3117,FA_out_3117}=FA_cout_2662+FA_out_2669+FA_cout_2713;
  assign {FA_cout_3118,FA_out_3118}=FA_cout_2663+FA_out_2684+FA_cout_2723;
  assign {FA_cout_3119,FA_out_3119}=FA_out_2665+FA_cout_2709+FA_out_2717;
  assign {FA_cout_3120,FA_out_3120}=FA_cout_2666+FA_out_2687+FA_cout_2742;
  assign {FA_cout_3121,FA_out_3121}=FA_out_2668+FA_cout_2736+FA_out_2744;
  assign {FA_cout_3122,FA_out_3122}=FA_cout_2669+FA_out_2690+FA_cout_2721;
  assign {FA_cout_3123,FA_out_3123}=FA_cout_2684+FA_out_2692+FA_cout_2731;
  assign {FA_cout_3124,FA_out_3124}=FA_out_2686+FA_cout_2717+FA_out_2725;
  assign {FA_cout_3125,FA_out_3125}=FA_cout_2687+FA_out_2695+FA_cout_2758;
  assign {FA_cout_3126,FA_out_3126}=FA_out_2689+FA_cout_2744+FA_out_2760;
  assign {FA_cout_3127,FA_out_3127}=FA_cout_2690+FA_out_2698+FA_cout_2729;
  assign {FA_cout_3128,FA_out_3128}=FA_out_2676+HA_cout_103+HA_out_104;
  assign {FA_cout_3129,FA_out_3129}=FA_out_2677+HA_cout_104+FA_out_2747;
  assign {FA_cout_3130,FA_out_3130}=FA_out_2678+FA_cout_2747+FA_out_2748;
  assign {FA_cout_3131,FA_out_3131}=FA_out_2679+FA_cout_2748+FA_out_2749;
  assign {FA_cout_3132,FA_out_3132}=FA_out_2680+FA_cout_2749+FA_out_2750;
  assign {FA_cout_3133,FA_out_3133}=FA_out_2681+FA_cout_2750+FA_out_2751;
  assign {FA_cout_3134,FA_out_3134}=FA_out_2682+FA_cout_2751+FA_out_2752;
  assign {FA_cout_3135,FA_out_3135}=FA_out_2683+FA_cout_2752+FA_out_2753;
  assign {FA_cout_3136,FA_out_3136}=FA_out_2691+FA_cout_2753+FA_out_2754;
  assign {FA_cout_3137,FA_out_3137}=FA_cout_2692+FA_out_2700+FA_cout_2739;
  assign {FA_cout_3138,FA_out_3138}=FA_out_2694+FA_cout_2725+FA_out_2733;
  assign {FA_cout_3139,FA_out_3139}=FA_cout_2695+FA_out_2703+FA_cout_2766;
  assign {FA_cout_3140,FA_out_3140}=FA_out_2697+FA_cout_2760+FA_out_2768;
  assign {FA_cout_3141,FA_out_3141}=FA_cout_2698+FA_out_2706+FA_cout_2737;
  assign {FA_cout_3142,FA_out_3142}=FA_out_2699+FA_cout_2754+FA_out_2771;
  assign {FA_cout_3143,FA_out_3143}=FA_cout_2700+FA_out_2708+FA_cout_2755;
  assign {FA_cout_3144,FA_out_3144}=FA_out_2702+FA_cout_2733+FA_out_2741;
  assign {FA_cout_3145,FA_out_3145}=FA_cout_2703+FA_out_2711+FA_cout_2775;
  assign {FA_cout_3146,FA_out_3146}=FA_out_2705+FA_cout_2768+FA_out_2777;
  assign {FA_cout_3147,FA_out_3147}=FA_cout_2706+FA_out_2714+FA_cout_2745;
  assign {FA_cout_3148,FA_out_3148}=FA_out_2707+FA_cout_2771+FA_out_2780;
  assign {FA_cout_3149,FA_out_3149}=FA_cout_2708+FA_out_2716+FA_cout_2763;
  assign {FA_cout_3150,FA_out_3150}=FA_out_2710+FA_cout_2741+FA_out_2757;
  assign {FA_cout_3151,FA_out_3151}=FA_cout_2711+FA_out_2719+FA_cout_2784;
  assign {FA_cout_3152,FA_out_3152}=FA_out_2713+FA_cout_2777+FA_out_2786;
  assign {FA_cout_3153,FA_out_3153}=FA_cout_2714+FA_out_2722+FA_cout_2761;
  assign {FA_cout_3154,FA_out_3154}=FA_out_2715+FA_cout_2780+FA_out_2789;
  assign {FA_cout_3155,FA_out_3155}=FA_cout_2716+FA_out_2724+FA_cout_2772;
  assign {FA_cout_3156,FA_out_3156}=FA_out_2718+FA_cout_2757+FA_out_2765;
  assign {FA_cout_3157,FA_out_3157}=FA_cout_2719+FA_out_2727+FA_cout_2790;
  assign {FA_cout_3158,FA_out_3158}=FA_out_2721+FA_cout_2786+HA_out_109;
  assign {FA_cout_3159,FA_out_3159}=FA_cout_2722+FA_out_2730+FA_cout_2769;
  assign {FA_cout_3160,FA_out_3160}=FA_out_2723+FA_cout_2789+HA_out_113;
  assign {FA_cout_3161,FA_out_3161}=FA_cout_2724+FA_out_2732+FA_cout_2781;
  assign {FA_cout_3162,FA_out_3162}=FA_out_2726+FA_cout_2765+FA_out_2774;
  assign {FA_cout_3163,FA_out_3163}=FA_cout_2727+FA_out_2735+HA_cout_116;
  assign {FA_cout_3164,FA_out_3164}=FA_out_2729+HA_cout_109+HA_out_118;
  assign {FA_cout_3165,FA_out_3165}=FA_cout_2730+FA_out_2738+FA_cout_2778;
  assign {FA_cout_3166,FA_out_3166}=FA_out_2731+HA_cout_113+HA_out_120;
  assign {FA_cout_3167,FA_out_3167}=FA_cout_2732+FA_out_2740+HA_cout_105;
  assign {FA_cout_3168,FA_out_3168}=FA_out_2734+FA_cout_2774+FA_out_2783;
  assign {FA_cout_3169,FA_out_3169}=FA_cout_2735+FA_out_2743+HA_cout_122;
  assign {FA_cout_3170,FA_out_3170}=FA_out_2737+HA_cout_118+HA_out_123;
  assign {FA_cout_3171,FA_out_3171}=FA_cout_2738+FA_out_2746+FA_cout_2787;
  assign {FA_cout_3172,FA_out_3172}=FA_out_2739+HA_cout_120+HA_out_125;
  assign {FA_cout_3173,FA_out_3173}=FA_cout_2740+FA_out_2756+HA_cout_114;
  assign {FA_cout_3174,FA_out_3174}=FA_out_2742+FA_cout_2783+HA_out_107;
  assign {FA_cout_3175,FA_out_3175}=FA_cout_2743+FA_out_2759+HA_cout_126;
  assign {FA_cout_3176,FA_out_3176}=FA_out_2745+HA_cout_123+REGS_1878;
  assign {FA_cout_3177,FA_out_3177}=FA_cout_2746+FA_out_2762+HA_cout_110;
  assign {FA_cout_3178,FA_out_3178}=FA_out_2755+HA_cout_125+REGS_1865;
  assign {FA_cout_3179,FA_out_3179}=FA_cout_2756+FA_out_2764+REGS_1846;
  assign {FA_cout_3180,FA_out_3180}=FA_out_2758+HA_cout_107+REGS_1798;
  assign {FA_cout_3181,FA_out_3181}=FA_cout_2762+FA_out_2770+REGS_1838;
  assign {FA_cout_3182,FA_out_3182}=FA_cout_2764+FA_out_2773+REGS_1867;
  assign {FA_cout_3183,FA_out_3183}=FA_cout_2770+FA_out_2779+REGS_1860;
  assign {FA_cout_3184,FA_out_3184}=FA_cout_2794+FA_out_2795+HA_out_88;
  assign {FA_cout_3185,FA_out_3185}=FA_cout_2795+FA_out_2796+HA_out_89;
  assign {FA_cout_3186,FA_out_3186}=FA_cout_2796+FA_out_2797+FA_out_2270;
  assign {FA_cout_3187,FA_out_3187}=FA_cout_2797+FA_out_2798+FA_out_2271;
  assign {FA_cout_3188,FA_out_3188}=FA_cout_2798+FA_out_2799+HA_out_131;
  assign {FA_cout_3189,FA_out_3189}=FA_cout_2799+FA_out_2800+HA_cout_131;
  assign {FA_cout_3190,FA_out_3190}=FA_cout_2800+FA_out_2801+HA_cout_132;
  assign {FA_cout_3191,FA_out_3191}=FA_cout_2801+FA_out_2802+HA_cout_133;
  assign {FA_cout_3192,FA_out_3192}=FA_cout_2802+FA_out_2803+FA_cout_2857;
  assign {FA_cout_3193,FA_out_3193}=FA_cout_2803+FA_out_2804+FA_cout_2858;
  assign {FA_cout_3194,FA_out_3194}=FA_cout_2804+FA_out_2805+FA_cout_2859;
  assign {FA_cout_3195,FA_out_3195}=FA_cout_2805+FA_out_2806+FA_cout_2860;
  assign {FA_cout_3196,FA_out_3196}=FA_cout_2806+FA_out_2807+FA_cout_2861;
  assign {FA_cout_3197,FA_out_3197}=FA_cout_2807+FA_out_2808+FA_cout_2862;
  assign {FA_cout_3198,FA_out_3198}=FA_cout_2808+FA_out_2809+FA_cout_2863;
  assign {FA_cout_3199,FA_out_3199}=FA_cout_2809+FA_out_2810+FA_cout_2864;
  assign {FA_cout_3200,FA_out_3200}=FA_cout_2810+FA_out_2811+FA_cout_2865;
  assign {FA_cout_3201,FA_out_3201}=FA_cout_2811+FA_out_2812+FA_cout_2866;
  assign {FA_cout_3202,FA_out_3202}=FA_cout_2812+FA_out_2813+FA_cout_2867;
  assign {FA_cout_3203,FA_out_3203}=FA_cout_2813+FA_out_2814+FA_cout_2868;
  assign {FA_cout_3204,FA_out_3204}=FA_cout_2814+FA_out_2815+FA_cout_2869;
  assign {FA_cout_3205,FA_out_3205}=FA_cout_2815+FA_out_2816+FA_cout_2870;
  assign {FA_cout_3206,FA_out_3206}=FA_cout_2816+FA_out_2817+FA_cout_2871;
  assign {FA_cout_3207,FA_out_3207}=FA_cout_2817+FA_out_2818+FA_cout_2872;
  assign {FA_cout_3208,FA_out_3208}=FA_cout_2818+FA_out_2819+FA_cout_2873;
  assign {FA_cout_3209,FA_out_3209}=FA_cout_2819+FA_out_2820+FA_cout_2874;
  assign {FA_cout_3210,FA_out_3210}=FA_cout_2820+FA_out_2821+FA_cout_2875;
  assign {FA_cout_3211,FA_out_3211}=FA_cout_2821+FA_out_2822+FA_cout_2876;
  assign {FA_cout_3212,FA_out_3212}=FA_cout_2822+FA_out_2823+FA_cout_2877;
  assign {FA_cout_3213,FA_out_3213}=FA_cout_2823+FA_out_2824+FA_cout_2878;
  assign {FA_cout_3214,FA_out_3214}=FA_cout_2824+FA_out_2825+FA_cout_2879;
  assign {FA_cout_3215,FA_out_3215}=FA_cout_2825+FA_out_2826+FA_cout_2880;
  assign {FA_cout_3216,FA_out_3216}=FA_cout_2826+FA_out_2827+FA_cout_2881;
  assign {FA_cout_3217,FA_out_3217}=FA_cout_2827+FA_out_2828+FA_cout_2882;
  assign {FA_cout_3218,FA_out_3218}=FA_cout_2828+FA_out_2829+FA_cout_2883;
  assign {FA_cout_3219,FA_out_3219}=FA_cout_2829+FA_out_2830+FA_cout_2884;
  assign {FA_cout_3220,FA_out_3220}=FA_cout_2830+FA_out_2831+FA_cout_2885;
  assign {FA_cout_3221,FA_out_3221}=FA_cout_2831+FA_out_2832+FA_cout_2886;
  assign {FA_cout_3222,FA_out_3222}=FA_cout_2832+FA_out_2833+FA_cout_2887;
  assign {FA_cout_3223,FA_out_3223}=FA_cout_2833+FA_out_2834+FA_cout_2888;
  assign {FA_cout_3224,FA_out_3224}=FA_cout_2834+FA_out_2835+FA_cout_2889;
  assign {FA_cout_3225,FA_out_3225}=FA_cout_2835+FA_out_2836+FA_cout_2890;
  assign {FA_cout_3226,FA_out_3226}=FA_cout_2836+FA_out_2837+FA_cout_2891;
  assign {FA_cout_3227,FA_out_3227}=FA_cout_2837+FA_out_2838+FA_cout_2892;
  assign {FA_cout_3228,FA_out_3228}=FA_cout_2838+FA_out_2839+FA_cout_2893;
  assign {FA_cout_3229,FA_out_3229}=FA_cout_2839+FA_out_2840+FA_cout_2894;
  assign {FA_cout_3230,FA_out_3230}=FA_cout_2840+FA_out_2841+FA_cout_2895;
  assign {FA_cout_3231,FA_out_3231}=FA_cout_2841+FA_out_2842+FA_cout_2896;
  assign {FA_cout_3232,FA_out_3232}=FA_cout_2842+FA_out_2843+FA_cout_2897;
  assign {FA_cout_3233,FA_out_3233}=FA_cout_2843+FA_out_2844+FA_cout_2898;
  assign {FA_cout_3234,FA_out_3234}=FA_cout_2844+FA_out_2845+FA_cout_2899;
  assign {FA_cout_3235,FA_out_3235}=FA_cout_2845+FA_out_2846+FA_cout_2900;
  assign {FA_cout_3236,FA_out_3236}=FA_cout_2846+FA_out_2847+FA_cout_2901;
  assign {FA_cout_3237,FA_out_3237}=FA_cout_2847+FA_out_2848+FA_cout_2902;
  assign {FA_cout_3238,FA_out_3238}=FA_cout_2848+FA_out_2849+FA_cout_2903;
  assign {FA_cout_3239,FA_out_3239}=FA_cout_2849+FA_out_2850+FA_cout_2904;
  assign {FA_cout_3240,FA_out_3240}=FA_cout_2850+FA_out_2851+FA_cout_2905;
  assign {FA_cout_3241,FA_out_3241}=FA_cout_2851+FA_out_2852+FA_cout_2906;
  assign {FA_cout_3242,FA_out_3242}=FA_cout_2852+FA_out_2853+FA_cout_2908;
  assign {FA_cout_3243,FA_out_3243}=FA_cout_2853+FA_out_2854+FA_cout_2910;
  assign {FA_cout_3244,FA_out_3244}=FA_cout_2854+FA_out_2855+FA_cout_2912;
  assign {FA_cout_3245,FA_out_3245}=FA_cout_2855+FA_out_2856+FA_cout_2914;
  assign {FA_cout_3246,FA_out_3246}=FA_cout_2856+FA_out_2907+FA_cout_2916;
  assign {FA_cout_3247,FA_out_3247}=FA_cout_2907+FA_out_2909+FA_cout_2918;
  assign {FA_cout_3248,FA_out_3248}=FA_out_2865+HA_cout_134+HA_out_135;
  assign {FA_cout_3249,FA_out_3249}=FA_out_2866+HA_cout_135+HA_out_136;
  assign {FA_cout_3250,FA_out_3250}=FA_out_2867+HA_cout_136+FA_out_2932;
  assign {FA_cout_3251,FA_out_3251}=FA_out_2868+FA_cout_2932+FA_out_2933;
  assign {FA_cout_3252,FA_out_3252}=FA_out_2869+FA_cout_2933+FA_out_2934;
  assign {FA_cout_3253,FA_out_3253}=FA_out_2870+FA_cout_2934+FA_out_2935;
  assign {FA_cout_3254,FA_out_3254}=FA_out_2871+FA_cout_2935+FA_out_2936;
  assign {FA_cout_3255,FA_out_3255}=FA_out_2872+FA_cout_2936+FA_out_2937;
  assign {FA_cout_3256,FA_out_3256}=FA_out_2873+FA_cout_2937+FA_out_2938;
  assign {FA_cout_3257,FA_out_3257}=FA_out_2874+FA_cout_2938+FA_out_2939;
  assign {FA_cout_3258,FA_out_3258}=FA_out_2875+FA_cout_2939+FA_out_2940;
  assign {FA_cout_3259,FA_out_3259}=FA_out_2876+FA_cout_2940+FA_out_2941;
  assign {FA_cout_3260,FA_out_3260}=FA_out_2877+FA_cout_2941+FA_out_2942;
  assign {FA_cout_3261,FA_out_3261}=FA_out_2878+FA_cout_2942+FA_out_2943;
  assign {FA_cout_3262,FA_out_3262}=FA_out_2879+FA_cout_2943+FA_out_2944;
  assign {FA_cout_3263,FA_out_3263}=FA_out_2880+FA_cout_2944+FA_out_2945;
  assign {FA_cout_3264,FA_out_3264}=FA_out_2881+FA_cout_2945+FA_out_2946;
  assign {FA_cout_3265,FA_out_3265}=FA_out_2882+FA_cout_2946+FA_out_2947;
  assign {FA_cout_3266,FA_out_3266}=FA_out_2883+FA_cout_2947+FA_out_2948;
  assign {FA_cout_3267,FA_out_3267}=FA_out_2884+FA_cout_2948+FA_out_2949;
  assign {FA_cout_3268,FA_out_3268}=FA_out_2885+FA_cout_2949+FA_out_2950;
  assign {FA_cout_3269,FA_out_3269}=FA_out_2886+FA_cout_2950+FA_out_2951;
  assign {FA_cout_3270,FA_out_3270}=FA_out_2887+FA_cout_2951+FA_out_2952;
  assign {FA_cout_3271,FA_out_3271}=FA_out_2888+FA_cout_2952+FA_out_2953;
  assign {FA_cout_3272,FA_out_3272}=FA_out_2889+FA_cout_2953+FA_out_2954;
  assign {FA_cout_3273,FA_out_3273}=FA_out_2890+FA_cout_2954+FA_out_2955;
  assign {FA_cout_3274,FA_out_3274}=FA_out_2891+FA_cout_2955+FA_out_2956;
  assign {FA_cout_3275,FA_out_3275}=FA_out_2892+FA_cout_2956+FA_out_2957;
  assign {FA_cout_3276,FA_out_3276}=FA_out_2893+FA_cout_2957+FA_out_2958;
  assign {FA_cout_3277,FA_out_3277}=FA_out_2894+FA_cout_2958+FA_out_2959;
  assign {FA_cout_3278,FA_out_3278}=FA_out_2895+FA_cout_2959+FA_out_2960;
  assign {FA_cout_3279,FA_out_3279}=FA_out_2896+FA_cout_2960+FA_out_2961;
  assign {FA_cout_3280,FA_out_3280}=FA_out_2897+FA_cout_2961+FA_out_2962;
  assign {FA_cout_3281,FA_out_3281}=FA_out_2898+FA_cout_2962+FA_out_2963;
  assign {FA_cout_3282,FA_out_3282}=FA_out_2899+FA_cout_2963+FA_out_2964;
  assign {FA_cout_3283,FA_out_3283}=FA_out_2900+FA_cout_2964+FA_out_2965;
  assign {FA_cout_3284,FA_out_3284}=FA_out_2901+FA_cout_2965+FA_out_2966;
  assign {FA_cout_3285,FA_out_3285}=FA_out_2902+FA_cout_2966+FA_out_2967;
  assign {FA_cout_3286,FA_out_3286}=FA_out_2903+FA_cout_2967+FA_out_2968;
  assign {FA_cout_3287,FA_out_3287}=FA_out_2904+FA_cout_2968+FA_out_2969;
  assign {FA_cout_3288,FA_out_3288}=FA_out_2905+FA_cout_2969+FA_out_2970;
  assign {FA_cout_3289,FA_out_3289}=FA_out_2906+FA_cout_2970+FA_out_2971;
  assign {FA_cout_3290,FA_out_3290}=FA_out_2908+FA_cout_2971+FA_out_2974;
  assign {FA_cout_3291,FA_out_3291}=FA_cout_2909+FA_out_2911+FA_cout_2920;
  assign {FA_cout_3292,FA_out_3292}=FA_out_2910+FA_cout_2974+FA_out_2977;
  assign {FA_cout_3293,FA_out_3293}=FA_cout_2911+FA_out_2913+FA_cout_2922;
  assign {FA_cout_3294,FA_out_3294}=FA_out_2912+FA_cout_2977+FA_out_2980;
  assign {FA_cout_3295,FA_out_3295}=FA_cout_2913+FA_out_2915+FA_cout_2924;
  assign {FA_cout_3296,FA_out_3296}=FA_out_2914+FA_cout_2980+FA_out_2983;
  assign {FA_cout_3297,FA_out_3297}=FA_cout_2915+FA_out_2917+FA_cout_2926;
  assign {FA_cout_3298,FA_out_3298}=FA_out_2916+FA_cout_2983+FA_out_2986;
  assign {FA_cout_3299,FA_out_3299}=FA_cout_2917+FA_out_2919+FA_cout_2928;
  assign {FA_cout_3300,FA_out_3300}=FA_out_2918+FA_cout_2986+FA_out_2989;
  assign {FA_cout_3301,FA_out_3301}=FA_cout_2919+FA_out_2921+FA_cout_2930;
  assign {FA_cout_3302,FA_out_3302}=FA_out_2920+FA_cout_2989+FA_out_2992;
  assign {FA_cout_3303,FA_out_3303}=FA_cout_2921+FA_out_2923+FA_cout_2972;
  assign {FA_cout_3304,FA_out_3304}=FA_out_2922+FA_cout_2992+FA_out_2995;
  assign {FA_cout_3305,FA_out_3305}=FA_cout_2923+FA_out_2925+FA_cout_2975;
  assign {FA_cout_3306,FA_out_3306}=FA_out_2924+FA_cout_2995+FA_out_3028;
  assign {FA_cout_3307,FA_out_3307}=FA_cout_2925+FA_out_2927+FA_cout_2978;
  assign {FA_cout_3308,FA_out_3308}=FA_out_2926+FA_cout_3028+FA_out_3032;
  assign {FA_cout_3309,FA_out_3309}=FA_cout_2927+FA_out_2929+FA_cout_2981;
  assign {FA_cout_3310,FA_out_3310}=FA_out_2928+FA_cout_3032+FA_out_3036;
  assign {FA_cout_3311,FA_out_3311}=FA_cout_2929+FA_out_2931+FA_cout_2984;
  assign {FA_cout_3312,FA_out_3312}=FA_out_2930+FA_cout_3036+FA_out_3040;
  assign {FA_cout_3313,FA_out_3313}=FA_cout_2931+FA_out_2973+FA_cout_2987;
  assign {FA_cout_3314,FA_out_3314}=FA_out_2972+FA_cout_3040+FA_out_3044;
  assign {FA_cout_3315,FA_out_3315}=FA_cout_2973+FA_out_2976+FA_cout_2990;
  assign {FA_cout_3316,FA_out_3316}=FA_out_2975+FA_cout_3044+FA_out_3048;
  assign {FA_cout_3317,FA_out_3317}=FA_cout_2976+FA_out_2979+FA_cout_2993;
  assign {FA_cout_3318,FA_out_3318}=FA_out_2978+FA_cout_3048+FA_out_3052;
  assign {FA_cout_3319,FA_out_3319}=FA_cout_2979+FA_out_2982+FA_cout_2996;
  assign {FA_cout_3320,FA_out_3320}=FA_out_2981+FA_cout_3052+FA_out_3056;
  assign {FA_cout_3321,FA_out_3321}=FA_cout_2982+FA_out_2985+FA_cout_3029;
  assign {FA_cout_3322,FA_out_3322}=FA_out_2984+FA_cout_3056+FA_out_3060;
  assign {FA_cout_3323,FA_out_3323}=FA_cout_2985+FA_out_2988+FA_cout_3033;
  assign {FA_cout_3324,FA_out_3324}=FA_out_2987+FA_cout_3060+FA_out_3064;
  assign {FA_cout_3325,FA_out_3325}=FA_cout_2988+FA_out_2991+FA_cout_3037;
  assign {FA_cout_3326,FA_out_3326}=FA_out_2990+FA_cout_3064+FA_out_3068;
  assign {FA_cout_3327,FA_out_3327}=FA_cout_2991+FA_out_2994+FA_cout_3041;
  assign {FA_cout_3328,FA_out_3328}=FA_out_2993+FA_cout_3068+FA_out_3072;
  assign {FA_cout_3329,FA_out_3329}=FA_cout_2994+FA_out_2997+FA_cout_3045;
  assign {FA_cout_3330,FA_out_3330}=FA_out_2996+FA_cout_3072+FA_out_3095;
  assign {FA_cout_3331,FA_out_3331}=FA_cout_2997+FA_out_3030+FA_cout_3049;
  assign {FA_cout_3332,FA_out_3332}=FA_cout_3001+FA_out_3002+REGS_1211;
  assign {FA_cout_3333,FA_out_3333}=FA_cout_3002+FA_out_3003+REGS_1212;
  assign {FA_cout_3334,FA_out_3334}=FA_cout_3003+FA_out_3004+HA_out_99;
  assign {FA_cout_3335,FA_out_3335}=FA_cout_3004+FA_out_3005+HA_out_141;
  assign {FA_cout_3336,FA_out_3336}=FA_cout_3005+FA_out_3006+HA_cout_141;
  assign {FA_cout_3337,FA_out_3337}=FA_cout_3006+FA_out_3007+HA_cout_142;
  assign {FA_cout_3338,FA_out_3338}=FA_cout_3007+FA_out_3008+HA_cout_143;
  assign {FA_cout_3339,FA_out_3339}=FA_cout_3008+FA_out_3009+HA_cout_144;
  assign {FA_cout_3340,FA_out_3340}=FA_cout_3009+FA_out_3010+FA_cout_3075;
  assign {FA_cout_3341,FA_out_3341}=FA_cout_3010+FA_out_3011+FA_cout_3076;
  assign {FA_cout_3342,FA_out_3342}=FA_cout_3011+FA_out_3012+FA_cout_3077;
  assign {FA_cout_3343,FA_out_3343}=FA_cout_3012+FA_out_3013+FA_cout_3078;
  assign {FA_cout_3344,FA_out_3344}=FA_cout_3013+FA_out_3014+FA_cout_3079;
  assign {FA_cout_3345,FA_out_3345}=FA_cout_3014+FA_out_3015+FA_cout_3080;
  assign {FA_cout_3346,FA_out_3346}=FA_cout_3015+FA_out_3016+FA_cout_3081;
  assign {FA_cout_3347,FA_out_3347}=FA_cout_3016+FA_out_3017+FA_cout_3082;
  assign {FA_cout_3348,FA_out_3348}=FA_cout_3017+FA_out_3018+FA_cout_3083;
  assign {FA_cout_3349,FA_out_3349}=FA_cout_3018+FA_out_3019+FA_cout_3084;
  assign {FA_cout_3350,FA_out_3350}=FA_cout_3019+FA_out_3020+FA_cout_3085;
  assign {FA_cout_3351,FA_out_3351}=FA_cout_3020+FA_out_3021+FA_cout_3086;
  assign {FA_cout_3352,FA_out_3352}=FA_cout_3021+FA_out_3022+FA_cout_3087;
  assign {FA_cout_3353,FA_out_3353}=FA_cout_3022+FA_out_3023+FA_cout_3088;
  assign {FA_cout_3354,FA_out_3354}=FA_cout_3023+FA_out_3024+FA_cout_3089;
  assign {FA_cout_3355,FA_out_3355}=FA_cout_3024+FA_out_3025+FA_cout_3090;
  assign {FA_cout_3356,FA_out_3356}=FA_cout_3025+FA_out_3026+FA_cout_3091;
  assign {FA_cout_3357,FA_out_3357}=FA_cout_3026+FA_out_3027+FA_cout_3092;
  assign {FA_cout_3358,FA_out_3358}=FA_cout_3027+FA_out_3031+FA_cout_3093;
  assign {FA_cout_3359,FA_out_3359}=FA_out_3029+FA_cout_3095+FA_out_3100;
  assign {FA_cout_3360,FA_out_3360}=FA_cout_3030+FA_out_3034+FA_cout_3053;
  assign {FA_cout_3361,FA_out_3361}=FA_cout_3031+FA_out_3035+FA_cout_3098;
  assign {FA_cout_3362,FA_out_3362}=FA_out_3033+FA_cout_3100+FA_out_3105;
  assign {FA_cout_3363,FA_out_3363}=FA_cout_3034+FA_out_3038+FA_cout_3057;
  assign {FA_cout_3364,FA_out_3364}=FA_cout_3035+FA_out_3039+FA_cout_3103;
  assign {FA_cout_3365,FA_out_3365}=FA_out_3037+FA_cout_3105+FA_out_3110;
  assign {FA_cout_3366,FA_out_3366}=FA_cout_3038+FA_out_3042+FA_cout_3061;
  assign {FA_cout_3367,FA_out_3367}=FA_cout_3039+FA_out_3043+FA_cout_3108;
  assign {FA_cout_3368,FA_out_3368}=FA_out_3041+FA_cout_3110+FA_out_3115;
  assign {FA_cout_3369,FA_out_3369}=FA_cout_3042+FA_out_3046+FA_cout_3065;
  assign {FA_cout_3370,FA_out_3370}=FA_cout_3043+FA_out_3047+FA_cout_3113;
  assign {FA_cout_3371,FA_out_3371}=FA_out_3045+FA_cout_3115+FA_out_3120;
  assign {FA_cout_3372,FA_out_3372}=FA_cout_3046+FA_out_3050+FA_cout_3069;
  assign {FA_cout_3373,FA_out_3373}=FA_cout_3047+FA_out_3051+FA_cout_3118;
  assign {FA_cout_3374,FA_out_3374}=FA_out_3049+FA_cout_3120+FA_out_3125;
  assign {FA_cout_3375,FA_out_3375}=FA_cout_3050+FA_out_3054+FA_cout_3073;
  assign {FA_cout_3376,FA_out_3376}=FA_cout_3051+FA_out_3055+FA_cout_3123;
  assign {FA_cout_3377,FA_out_3377}=FA_out_3053+FA_cout_3125+FA_out_3139;
  assign {FA_cout_3378,FA_out_3378}=FA_cout_3054+FA_out_3058+FA_cout_3096;
  assign {FA_cout_3379,FA_out_3379}=FA_cout_3055+FA_out_3059+FA_cout_3137;
  assign {FA_cout_3380,FA_out_3380}=FA_out_3057+FA_cout_3139+FA_out_3145;
  assign {FA_cout_3381,FA_out_3381}=FA_cout_3058+FA_out_3062+FA_cout_3101;
  assign {FA_cout_3382,FA_out_3382}=FA_cout_3059+FA_out_3063+FA_cout_3143;
  assign {FA_cout_3383,FA_out_3383}=FA_out_3061+FA_cout_3145+FA_out_3151;
  assign {FA_cout_3384,FA_out_3384}=FA_cout_3062+FA_out_3066+FA_cout_3106;
  assign {FA_cout_3385,FA_out_3385}=FA_cout_3063+FA_out_3067+FA_cout_3149;
  assign {FA_cout_3386,FA_out_3386}=FA_out_3065+FA_cout_3151+FA_out_3157;
  assign {FA_cout_3387,FA_out_3387}=FA_cout_3066+FA_out_3070+FA_cout_3111;
  assign {FA_cout_3388,FA_out_3388}=FA_cout_3067+FA_out_3071+FA_cout_3155;
  assign {FA_cout_3389,FA_out_3389}=FA_out_3069+FA_cout_3157+FA_out_3163;
  assign {FA_cout_3390,FA_out_3390}=FA_cout_3070+FA_out_3074+FA_cout_3116;
  assign {FA_cout_3391,FA_out_3391}=FA_cout_3071+FA_out_3094+FA_cout_3161;
  assign {FA_cout_3392,FA_out_3392}=FA_out_3073+FA_cout_3163+FA_out_3169;
  assign {FA_cout_3393,FA_out_3393}=FA_cout_3074+FA_out_3097+FA_cout_3121;
  assign {FA_cout_3394,FA_out_3394}=FA_cout_3094+FA_out_3099+FA_cout_3167;
  assign {FA_cout_3395,FA_out_3395}=FA_out_3096+FA_cout_3169+FA_out_3175;
  assign {FA_cout_3396,FA_out_3396}=FA_cout_3097+FA_out_3102+FA_cout_3126;
  assign {FA_cout_3397,FA_out_3397}=FA_out_3082+HA_cout_145+HA_out_146;
  assign {FA_cout_3398,FA_out_3398}=FA_out_3083+HA_cout_146+HA_out_147;
  assign {FA_cout_3399,FA_out_3399}=FA_out_3084+HA_cout_147+HA_out_148;
  assign {FA_cout_3400,FA_out_3400}=FA_out_3085+HA_cout_148+FA_out_3128;
  assign {FA_cout_3401,FA_out_3401}=FA_out_3086+FA_cout_3128+FA_out_3129;
  assign {FA_cout_3402,FA_out_3402}=FA_out_3087+FA_cout_3129+FA_out_3130;
  assign {FA_cout_3403,FA_out_3403}=FA_out_3088+FA_cout_3130+FA_out_3131;
  assign {FA_cout_3404,FA_out_3404}=FA_out_3089+FA_cout_3131+FA_out_3132;
  assign {FA_cout_3405,FA_out_3405}=FA_out_3090+FA_cout_3132+FA_out_3133;
  assign {FA_cout_3406,FA_out_3406}=FA_out_3091+FA_cout_3133+FA_out_3134;
  assign {FA_cout_3407,FA_out_3407}=FA_out_3092+FA_cout_3134+FA_out_3135;
  assign {FA_cout_3408,FA_out_3408}=FA_out_3093+FA_cout_3135+FA_out_3136;
  assign {FA_cout_3409,FA_out_3409}=FA_out_3098+FA_cout_3136+FA_out_3142;
  assign {FA_cout_3410,FA_out_3410}=FA_cout_3099+FA_out_3104+FA_cout_3173;
  assign {FA_cout_3411,FA_out_3411}=FA_out_3101+FA_cout_3175+HA_out_149;
  assign {FA_cout_3412,FA_out_3412}=FA_cout_3102+FA_out_3107+FA_cout_3140;
  assign {FA_cout_3413,FA_out_3413}=FA_out_3103+FA_cout_3142+FA_out_3148;
  assign {FA_cout_3414,FA_out_3414}=FA_cout_3104+FA_out_3109+FA_cout_3179;
  assign {FA_cout_3415,FA_out_3415}=FA_out_3106+HA_cout_149+HA_out_152;
  assign {FA_cout_3416,FA_out_3416}=FA_cout_3107+FA_out_3112+FA_cout_3146;
  assign {FA_cout_3417,FA_out_3417}=FA_out_3108+FA_cout_3148+FA_out_3154;
  assign {FA_cout_3418,FA_out_3418}=FA_cout_3109+FA_out_3114+FA_cout_3182;
  assign {FA_cout_3419,FA_out_3419}=FA_out_3111+HA_cout_152+HA_out_155;
  assign {FA_cout_3420,FA_out_3420}=FA_cout_3112+FA_out_3117+FA_cout_3152;
  assign {FA_cout_3421,FA_out_3421}=FA_out_3113+FA_cout_3154+FA_out_3160;
  assign {FA_cout_3422,FA_out_3422}=FA_cout_3114+FA_out_3119+HA_cout_153;
  assign {FA_cout_3423,FA_out_3423}=FA_out_3116+HA_cout_155+HA_out_158;
  assign {FA_cout_3424,FA_out_3424}=FA_cout_3117+FA_out_3122+FA_cout_3158;
  assign {FA_cout_3425,FA_out_3425}=FA_out_3118+FA_cout_3160+FA_out_3166;
  assign {FA_cout_3426,FA_out_3426}=FA_cout_3119+FA_out_3124+HA_cout_157;
  assign {FA_cout_3427,FA_out_3427}=FA_out_3121+HA_cout_158+HA_out_161;
  assign {FA_cout_3428,FA_out_3428}=FA_cout_3122+FA_out_3127+FA_cout_3164;
  assign {FA_cout_3429,FA_out_3429}=FA_out_3123+FA_cout_3166+FA_out_3172;
  assign {FA_cout_3430,FA_out_3430}=FA_cout_3124+FA_out_3138+HA_cout_160;
  assign {FA_cout_3431,FA_out_3431}=FA_out_3126+HA_cout_161+HA_out_166;
  assign {FA_cout_3432,FA_out_3432}=FA_cout_3127+FA_out_3141+FA_cout_3170;
  assign {FA_cout_3433,FA_out_3433}=FA_out_3137+FA_cout_3172+FA_out_3178;
  assign {FA_cout_3434,FA_out_3434}=FA_cout_3138+FA_out_3144+HA_cout_165;
  assign {FA_cout_3435,FA_out_3435}=FA_out_3140+HA_cout_166+REGS_1855;
  assign {FA_cout_3436,FA_out_3436}=FA_cout_3141+FA_out_3147+FA_cout_3176;
  assign {FA_cout_3437,FA_out_3437}=FA_out_3143+FA_cout_3178+FA_out_2763;
  assign {FA_cout_3438,FA_out_3438}=FA_cout_3144+FA_out_3150+HA_cout_168;
  assign {FA_cout_3439,FA_out_3439}=FA_cout_3147+FA_out_3153+HA_cout_150;
  assign {FA_cout_3440,FA_out_3440}=FA_cout_3153+FA_out_3159+FA_out_2778;
  assign {FA_cout_3441,FA_out_3441}=FA_cout_3159+FA_out_3165+FA_out_2787;
  assign {FA_cout_3442,FA_out_3442}=FA_cout_3165+FA_out_3171+HA_out_110;
  assign {FA_cout_3443,FA_out_3443}=FA_cout_3171+FA_out_3177+REGS_1810;
  assign {FA_cout_3444,FA_out_3444}=FA_cout_3188+FA_out_3189+HA_out_132;
  assign {FA_cout_3445,FA_out_3445}=FA_cout_3189+FA_out_3190+HA_out_133;
  assign {FA_cout_3446,FA_out_3446}=FA_cout_3190+FA_out_3191+FA_out_2857;
  assign {FA_cout_3447,FA_out_3447}=FA_cout_3191+FA_out_3192+FA_out_2858;
  assign {FA_cout_3448,FA_out_3448}=FA_cout_3192+FA_out_3193+FA_out_2859;
  assign {FA_cout_3449,FA_out_3449}=FA_cout_3193+FA_out_3194+FA_out_2860;
  assign {FA_cout_3450,FA_out_3450}=FA_cout_3194+FA_out_3195+HA_out_176;
  assign {FA_cout_3451,FA_out_3451}=FA_cout_3195+FA_out_3196+HA_cout_176;
  assign {FA_cout_3452,FA_out_3452}=FA_cout_3196+FA_out_3197+HA_cout_177;
  assign {FA_cout_3453,FA_out_3453}=FA_cout_3197+FA_out_3198+HA_cout_178;
  assign {FA_cout_3454,FA_out_3454}=FA_cout_3198+FA_out_3199+HA_cout_179;
  assign {FA_cout_3455,FA_out_3455}=FA_cout_3199+FA_out_3200+FA_cout_3248;
  assign {FA_cout_3456,FA_out_3456}=FA_cout_3200+FA_out_3201+FA_cout_3249;
  assign {FA_cout_3457,FA_out_3457}=FA_cout_3201+FA_out_3202+FA_cout_3250;
  assign {FA_cout_3458,FA_out_3458}=FA_cout_3202+FA_out_3203+FA_cout_3251;
  assign {FA_cout_3459,FA_out_3459}=FA_cout_3203+FA_out_3204+FA_cout_3252;
  assign {FA_cout_3460,FA_out_3460}=FA_cout_3204+FA_out_3205+FA_cout_3253;
  assign {FA_cout_3461,FA_out_3461}=FA_cout_3205+FA_out_3206+FA_cout_3254;
  assign {FA_cout_3462,FA_out_3462}=FA_cout_3206+FA_out_3207+FA_cout_3255;
  assign {FA_cout_3463,FA_out_3463}=FA_cout_3207+FA_out_3208+FA_cout_3256;
  assign {FA_cout_3464,FA_out_3464}=FA_cout_3208+FA_out_3209+FA_cout_3257;
  assign {FA_cout_3465,FA_out_3465}=FA_cout_3209+FA_out_3210+FA_cout_3258;
  assign {FA_cout_3466,FA_out_3466}=FA_cout_3210+FA_out_3211+FA_cout_3259;
  assign {FA_cout_3467,FA_out_3467}=FA_cout_3211+FA_out_3212+FA_cout_3260;
  assign {FA_cout_3468,FA_out_3468}=FA_cout_3212+FA_out_3213+FA_cout_3261;
  assign {FA_cout_3469,FA_out_3469}=FA_cout_3213+FA_out_3214+FA_cout_3262;
  assign {FA_cout_3470,FA_out_3470}=FA_cout_3214+FA_out_3215+FA_cout_3263;
  assign {FA_cout_3471,FA_out_3471}=FA_cout_3215+FA_out_3216+FA_cout_3264;
  assign {FA_cout_3472,FA_out_3472}=FA_cout_3216+FA_out_3217+FA_cout_3265;
  assign {FA_cout_3473,FA_out_3473}=FA_cout_3217+FA_out_3218+FA_cout_3266;
  assign {FA_cout_3474,FA_out_3474}=FA_cout_3218+FA_out_3219+FA_cout_3267;
  assign {FA_cout_3475,FA_out_3475}=FA_cout_3219+FA_out_3220+FA_cout_3268;
  assign {FA_cout_3476,FA_out_3476}=FA_cout_3220+FA_out_3221+FA_cout_3269;
  assign {FA_cout_3477,FA_out_3477}=FA_cout_3221+FA_out_3222+FA_cout_3270;
  assign {FA_cout_3478,FA_out_3478}=FA_cout_3222+FA_out_3223+FA_cout_3271;
  assign {FA_cout_3479,FA_out_3479}=FA_cout_3223+FA_out_3224+FA_cout_3272;
  assign {FA_cout_3480,FA_out_3480}=FA_cout_3224+FA_out_3225+FA_cout_3273;
  assign {FA_cout_3481,FA_out_3481}=FA_cout_3225+FA_out_3226+FA_cout_3274;
  assign {FA_cout_3482,FA_out_3482}=FA_cout_3226+FA_out_3227+FA_cout_3275;
  assign {FA_cout_3483,FA_out_3483}=FA_cout_3227+FA_out_3228+FA_cout_3276;
  assign {FA_cout_3484,FA_out_3484}=FA_cout_3228+FA_out_3229+FA_cout_3277;
  assign {FA_cout_3485,FA_out_3485}=FA_cout_3229+FA_out_3230+FA_cout_3278;
  assign {FA_cout_3486,FA_out_3486}=FA_cout_3230+FA_out_3231+FA_cout_3279;
  assign {FA_cout_3487,FA_out_3487}=FA_cout_3231+FA_out_3232+FA_cout_3280;
  assign {FA_cout_3488,FA_out_3488}=FA_cout_3232+FA_out_3233+FA_cout_3281;
  assign {FA_cout_3489,FA_out_3489}=FA_cout_3233+FA_out_3234+FA_cout_3282;
  assign {FA_cout_3490,FA_out_3490}=FA_cout_3234+FA_out_3235+FA_cout_3283;
  assign {FA_cout_3491,FA_out_3491}=FA_cout_3235+FA_out_3236+FA_cout_3284;
  assign {FA_cout_3492,FA_out_3492}=FA_cout_3236+FA_out_3237+FA_cout_3285;
  assign {FA_cout_3493,FA_out_3493}=FA_cout_3237+FA_out_3238+FA_cout_3286;
  assign {FA_cout_3494,FA_out_3494}=FA_cout_3238+FA_out_3239+FA_cout_3287;
  assign {FA_cout_3495,FA_out_3495}=FA_cout_3239+FA_out_3240+FA_cout_3288;
  assign {FA_cout_3496,FA_out_3496}=FA_cout_3240+FA_out_3241+FA_cout_3289;
  assign {FA_cout_3497,FA_out_3497}=FA_cout_3241+FA_out_3242+FA_cout_3290;
  assign {FA_cout_3498,FA_out_3498}=FA_cout_3242+FA_out_3243+FA_cout_3292;
  assign {FA_cout_3499,FA_out_3499}=FA_cout_3243+FA_out_3244+FA_cout_3294;
  assign {FA_cout_3500,FA_out_3500}=FA_cout_3244+FA_out_3245+FA_cout_3296;
  assign {FA_cout_3501,FA_out_3501}=FA_cout_3245+FA_out_3246+FA_cout_3298;
  assign {FA_cout_3502,FA_out_3502}=FA_cout_3246+FA_out_3247+FA_cout_3300;
  assign {FA_cout_3503,FA_out_3503}=FA_cout_3247+FA_out_3291+FA_cout_3302;
  assign {FA_cout_3504,FA_out_3504}=FA_cout_3291+FA_out_3293+FA_cout_3304;
  assign {FA_cout_3505,FA_out_3505}=FA_out_3258+HA_cout_180+HA_out_181;
  assign {FA_cout_3506,FA_out_3506}=FA_out_3259+HA_cout_181+HA_out_182;
  assign {FA_cout_3507,FA_out_3507}=FA_out_3260+HA_cout_182+HA_out_183;
  assign {FA_cout_3508,FA_out_3508}=FA_out_3261+HA_cout_183+HA_out_184;
  assign {FA_cout_3509,FA_out_3509}=FA_out_3262+HA_cout_184+HA_out_185;
  assign {FA_cout_3510,FA_out_3510}=FA_out_3263+HA_cout_185+HA_out_186;
  assign {FA_cout_3511,FA_out_3511}=FA_out_3264+HA_cout_186+FA_out_3332;
  assign {FA_cout_3512,FA_out_3512}=FA_out_3265+FA_cout_3332+FA_out_3333;
  assign {FA_cout_3513,FA_out_3513}=FA_out_3266+FA_cout_3333+FA_out_3334;
  assign {FA_cout_3514,FA_out_3514}=FA_out_3267+FA_cout_3334+FA_out_3335;
  assign {FA_cout_3515,FA_out_3515}=FA_out_3268+FA_cout_3335+FA_out_3336;
  assign {FA_cout_3516,FA_out_3516}=FA_out_3269+FA_cout_3336+FA_out_3337;
  assign {FA_cout_3517,FA_out_3517}=FA_out_3270+FA_cout_3337+FA_out_3338;
  assign {FA_cout_3518,FA_out_3518}=FA_out_3271+FA_cout_3338+FA_out_3339;
  assign {FA_cout_3519,FA_out_3519}=FA_out_3272+FA_cout_3339+FA_out_3340;
  assign {FA_cout_3520,FA_out_3520}=FA_out_3273+FA_cout_3340+FA_out_3341;
  assign {FA_cout_3521,FA_out_3521}=FA_out_3274+FA_cout_3341+FA_out_3342;
  assign {FA_cout_3522,FA_out_3522}=FA_out_3275+FA_cout_3342+FA_out_3343;
  assign {FA_cout_3523,FA_out_3523}=FA_out_3276+FA_cout_3343+FA_out_3344;
  assign {FA_cout_3524,FA_out_3524}=FA_out_3277+FA_cout_3344+FA_out_3345;
  assign {FA_cout_3525,FA_out_3525}=FA_out_3278+FA_cout_3345+FA_out_3346;
  assign {FA_cout_3526,FA_out_3526}=FA_out_3279+FA_cout_3346+FA_out_3347;
  assign {FA_cout_3527,FA_out_3527}=FA_out_3280+FA_cout_3347+FA_out_3348;
  assign {FA_cout_3528,FA_out_3528}=FA_out_3281+FA_cout_3348+FA_out_3349;
  assign {FA_cout_3529,FA_out_3529}=FA_out_3282+FA_cout_3349+FA_out_3350;
  assign {FA_cout_3530,FA_out_3530}=FA_out_3283+FA_cout_3350+FA_out_3351;
  assign {FA_cout_3531,FA_out_3531}=FA_out_3284+FA_cout_3351+FA_out_3352;
  assign {FA_cout_3532,FA_out_3532}=FA_out_3285+FA_cout_3352+FA_out_3353;
  assign {FA_cout_3533,FA_out_3533}=FA_out_3286+FA_cout_3353+FA_out_3354;
  assign {FA_cout_3534,FA_out_3534}=FA_out_3287+FA_cout_3354+FA_out_3355;
  assign {FA_cout_3535,FA_out_3535}=FA_out_3288+FA_cout_3355+FA_out_3356;
  assign {FA_cout_3536,FA_out_3536}=FA_out_3289+FA_cout_3356+FA_out_3357;
  assign {FA_cout_3537,FA_out_3537}=FA_out_3290+FA_cout_3357+FA_out_3358;
  assign {FA_cout_3538,FA_out_3538}=FA_out_3292+FA_cout_3358+FA_out_3361;
  assign {FA_cout_3539,FA_out_3539}=FA_cout_3293+FA_out_3295+FA_cout_3306;
  assign {FA_cout_3540,FA_out_3540}=FA_out_3294+FA_cout_3361+FA_out_3364;
  assign {FA_cout_3541,FA_out_3541}=FA_cout_3295+FA_out_3297+FA_cout_3308;
  assign {FA_cout_3542,FA_out_3542}=FA_out_3296+FA_cout_3364+FA_out_3367;
  assign {FA_cout_3543,FA_out_3543}=FA_cout_3297+FA_out_3299+FA_cout_3310;
  assign {FA_cout_3544,FA_out_3544}=FA_out_3298+FA_cout_3367+FA_out_3370;
  assign {FA_cout_3545,FA_out_3545}=FA_cout_3299+FA_out_3301+FA_cout_3312;
  assign {FA_cout_3546,FA_out_3546}=FA_out_3300+FA_cout_3370+FA_out_3373;
  assign {FA_cout_3547,FA_out_3547}=FA_cout_3301+FA_out_3303+FA_cout_3314;
  assign {FA_cout_3548,FA_out_3548}=FA_out_3302+FA_cout_3373+FA_out_3376;
  assign {FA_cout_3549,FA_out_3549}=FA_cout_3303+FA_out_3305+FA_cout_3316;
  assign {FA_cout_3550,FA_out_3550}=FA_out_3304+FA_cout_3376+FA_out_3379;
  assign {FA_cout_3551,FA_out_3551}=FA_cout_3305+FA_out_3307+FA_cout_3318;
  assign {FA_cout_3552,FA_out_3552}=FA_out_3306+FA_cout_3379+FA_out_3382;
  assign {FA_cout_3553,FA_out_3553}=FA_cout_3307+FA_out_3309+FA_cout_3320;
  assign {FA_cout_3554,FA_out_3554}=FA_out_3308+FA_cout_3382+FA_out_3385;
  assign {FA_cout_3555,FA_out_3555}=FA_cout_3309+FA_out_3311+FA_cout_3322;
  assign {FA_cout_3556,FA_out_3556}=FA_out_3310+FA_cout_3385+FA_out_3388;
  assign {FA_cout_3557,FA_out_3557}=FA_cout_3311+FA_out_3313+FA_cout_3324;
  assign {FA_cout_3558,FA_out_3558}=FA_out_3312+FA_cout_3388+FA_out_3391;
  assign {FA_cout_3559,FA_out_3559}=FA_cout_3313+FA_out_3315+FA_cout_3326;
  assign {FA_cout_3560,FA_out_3560}=FA_out_3314+FA_cout_3391+FA_out_3394;
  assign {FA_cout_3561,FA_out_3561}=FA_cout_3315+FA_out_3317+FA_cout_3328;
  assign {FA_cout_3562,FA_out_3562}=FA_out_3316+FA_cout_3394+FA_out_3410;
  assign {FA_cout_3563,FA_out_3563}=FA_cout_3317+FA_out_3319+FA_cout_3330;
  assign {FA_cout_3564,FA_out_3564}=FA_out_3318+FA_cout_3410+FA_out_3414;
  assign {FA_cout_3565,FA_out_3565}=FA_cout_3319+FA_out_3321+FA_cout_3359;
  assign {FA_cout_3566,FA_out_3566}=FA_out_3320+FA_cout_3414+FA_out_3418;
  assign {FA_cout_3567,FA_out_3567}=FA_cout_3321+FA_out_3323+FA_cout_3362;
  assign {FA_cout_3568,FA_out_3568}=FA_out_3322+FA_cout_3418+FA_out_3422;
  assign {FA_cout_3569,FA_out_3569}=FA_cout_3323+FA_out_3325+FA_cout_3365;
  assign {FA_cout_3570,FA_out_3570}=FA_out_3324+FA_cout_3422+FA_out_3426;
  assign {FA_cout_3571,FA_out_3571}=FA_cout_3325+FA_out_3327+FA_cout_3368;
  assign {FA_cout_3572,FA_out_3572}=FA_out_3326+FA_cout_3426+FA_out_3430;
  assign {FA_cout_3573,FA_out_3573}=FA_cout_3327+FA_out_3329+FA_cout_3371;
  assign {FA_cout_3574,FA_out_3574}=FA_out_3328+FA_cout_3430+FA_out_3434;
  assign {FA_cout_3575,FA_out_3575}=FA_cout_3329+FA_out_3331+FA_cout_3374;
  assign {FA_cout_3576,FA_out_3576}=FA_out_3330+FA_cout_3434+FA_out_3438;
  assign {FA_cout_3577,FA_out_3577}=FA_cout_3331+FA_out_3360+FA_cout_3377;
  assign {FA_cout_3578,FA_out_3578}=FA_out_3359+FA_cout_3438+HA_out_193;
  assign {FA_cout_3579,FA_out_3579}=FA_cout_3360+FA_out_3363+FA_cout_3380;
  assign {FA_cout_3580,FA_out_3580}=FA_out_3362+HA_cout_193+HA_out_195;
  assign {FA_cout_3581,FA_out_3581}=FA_cout_3363+FA_out_3366+FA_cout_3383;
  assign {FA_cout_3582,FA_out_3582}=FA_out_3365+HA_cout_195+HA_out_197;
  assign {FA_cout_3583,FA_out_3583}=FA_cout_3366+FA_out_3369+FA_cout_3386;
  assign {FA_cout_3584,FA_out_3584}=FA_out_3368+HA_cout_197+HA_out_199;
  assign {FA_cout_3585,FA_out_3585}=FA_cout_3369+FA_out_3372+FA_cout_3389;
  assign {FA_cout_3586,FA_out_3586}=FA_out_3371+HA_cout_199+HA_out_201;
  assign {FA_cout_3587,FA_out_3587}=FA_cout_3372+FA_out_3375+FA_cout_3392;
  assign {FA_cout_3588,FA_out_3588}=FA_out_3374+HA_cout_201+HA_out_203;
  assign {FA_cout_3589,FA_out_3589}=FA_cout_3375+FA_out_3378+FA_cout_3395;
  assign {FA_cout_3590,FA_out_3590}=FA_out_3377+HA_cout_203+HA_out_205;
  assign {FA_cout_3591,FA_out_3591}=FA_cout_3378+FA_out_3381+FA_cout_3411;
  assign {FA_cout_3592,FA_out_3592}=FA_out_3380+HA_cout_205+HA_out_207;
  assign {FA_cout_3593,FA_out_3593}=FA_cout_3381+FA_out_3384+FA_cout_3415;
  assign {FA_cout_3594,FA_out_3594}=FA_out_3383+HA_cout_207+FA_out_2790;
  assign {FA_cout_3595,FA_out_3595}=FA_cout_3384+FA_out_3387+FA_cout_3419;
  assign {FA_cout_3596,FA_out_3596}=FA_cout_3387+FA_out_3390+FA_cout_3423;
  assign {FA_cout_3597,FA_out_3597}=FA_cout_3390+FA_out_3393+FA_cout_3427;
  assign {FA_cout_3598,FA_out_3598}=FA_cout_3393+FA_out_3396+FA_cout_3431;
  assign {FA_cout_3599,FA_out_3599}=FA_cout_3396+FA_out_3412+FA_cout_3435;
  assign {FA_cout_3600,FA_out_3600}=FA_cout_3402+FA_out_3403+REGS_1782;
  assign {FA_cout_3601,FA_out_3601}=FA_cout_3403+FA_out_3404+REGS_1783;
  assign {FA_cout_3602,FA_out_3602}=FA_cout_3404+FA_out_3405+HA_out_111;
  assign {FA_cout_3603,FA_out_3603}=FA_cout_3405+FA_out_3406+HA_out_163;
  assign {FA_cout_3604,FA_out_3604}=FA_cout_3406+FA_out_3407+HA_out_211;
  assign {FA_cout_3605,FA_out_3605}=FA_cout_3407+FA_out_3408+HA_cout_211;
  assign {FA_cout_3606,FA_out_3606}=FA_cout_3408+FA_out_3409+HA_cout_212;
  assign {FA_cout_3607,FA_out_3607}=FA_cout_3412+FA_out_3416+HA_cout_191;
  assign {FA_cout_3608,FA_out_3608}=FA_cout_3416+FA_out_3420+FA_out_3158;
  assign {FA_cout_3609,FA_out_3609}=FA_cout_3420+FA_out_3424+FA_out_3164;
  assign {FA_cout_3610,FA_out_3610}=FA_cout_3424+FA_out_3428+FA_out_3170;
  assign {FA_cout_3611,FA_out_3611}=FA_cout_3428+FA_out_3432+FA_out_3176;
  assign {FA_cout_3612,FA_out_3612}=FA_cout_3432+FA_out_3436+HA_out_150;
  assign {FA_cout_3613,FA_out_3613}=FA_cout_3436+FA_out_3439+FA_out_2769;
  assign {FA_cout_3614,FA_out_3614}=REGS_1915+REGS_1979+REGS_2039;
  assign {FA_cout_3615,FA_out_3615}=REGS_1916+REGS_1980+REGS_2040;
  assign {FA_cout_3616,FA_out_3616}=REGS_1917+REGS_1981+REGS_2041;
  assign {FA_cout_3617,FA_out_3617}=REGS_1918+REGS_1982+REGS_2042;
  assign {FA_cout_3618,FA_out_3618}=REGS_1919+REGS_1983+REGS_2043;
  assign {FA_cout_3619,FA_out_3619}=REGS_1920+REGS_1984+REGS_2044;
  assign {FA_cout_3620,FA_out_3620}=REGS_1921+REGS_1985+REGS_2045;
  assign {FA_cout_3621,FA_out_3621}=REGS_1922+REGS_1986+REGS_2046;
  assign {FA_cout_3622,FA_out_3622}=REGS_1923+REGS_1987+REGS_2047;
  assign {FA_cout_3623,FA_out_3623}=REGS_1924+REGS_1988+REGS_2048;
  assign {FA_cout_3624,FA_out_3624}=REGS_1925+REGS_1989+REGS_2049;
  assign {FA_cout_3625,FA_out_3625}=REGS_1926+REGS_1990+REGS_2050;
  assign {FA_cout_3626,FA_out_3626}=REGS_1927+REGS_1991+REGS_2051;
  assign {FA_cout_3627,FA_out_3627}=REGS_1928+REGS_1992+REGS_2052;
  assign {FA_cout_3628,FA_out_3628}=REGS_1929+REGS_1993+REGS_2053;
  assign {FA_cout_3629,FA_out_3629}=REGS_1930+REGS_1994+REGS_2054;
  assign {FA_cout_3630,FA_out_3630}=REGS_1931+REGS_1995+REGS_2055;
  assign {FA_cout_3631,FA_out_3631}=REGS_1932+REGS_1996+REGS_2056;
  assign {FA_cout_3632,FA_out_3632}=REGS_1933+REGS_1997+REGS_2057;
  assign {FA_cout_3633,FA_out_3633}=REGS_1934+REGS_1998+REGS_2058;
  assign {FA_cout_3634,FA_out_3634}=REGS_1935+REGS_1999+REGS_2059;
  assign {FA_cout_3635,FA_out_3635}=REGS_1936+REGS_2000+REGS_2060;
  assign {FA_cout_3636,FA_out_3636}=REGS_1937+REGS_2001+REGS_2061;
  assign {FA_cout_3637,FA_out_3637}=REGS_1938+REGS_2002+REGS_2062;
  assign {FA_cout_3638,FA_out_3638}=REGS_1939+REGS_2003+REGS_2063;
  assign {FA_cout_3639,FA_out_3639}=REGS_1940+REGS_2004+REGS_2064;
  assign {FA_cout_3640,FA_out_3640}=REGS_1941+REGS_2005+REGS_2065;
  assign {FA_cout_3641,FA_out_3641}=REGS_1942+REGS_2006+REGS_2066;
  assign {FA_cout_3642,FA_out_3642}=REGS_1943+REGS_2007+REGS_2067;
  assign {FA_cout_3643,FA_out_3643}=REGS_1944+REGS_2008+REGS_2068;
  assign {FA_cout_3644,FA_out_3644}=REGS_1945+REGS_2009+REGS_2069;
  assign {FA_cout_3645,FA_out_3645}=REGS_1946+REGS_2010+REGS_2070;
  assign {FA_cout_3646,FA_out_3646}=REGS_1947+REGS_2011+REGS_2071;
  assign {FA_cout_3647,FA_out_3647}=REGS_1948+REGS_2012+REGS_2072;
  assign {FA_cout_3648,FA_out_3648}=REGS_1949+REGS_2013+REGS_2073;
  assign {FA_cout_3649,FA_out_3649}=REGS_1950+REGS_2014+REGS_2074;
  assign {FA_cout_3650,FA_out_3650}=REGS_1951+REGS_2015+REGS_2075;
  assign {FA_cout_3651,FA_out_3651}=REGS_1952+REGS_2016+REGS_2076;
  assign {FA_cout_3652,FA_out_3652}=REGS_1953+REGS_2017+REGS_2077;
  assign {FA_cout_3653,FA_out_3653}=REGS_1954+REGS_2018+REGS_2078;
  assign {FA_cout_3654,FA_out_3654}=REGS_1955+REGS_2019+REGS_2079;
  assign {FA_cout_3655,FA_out_3655}=REGS_1956+REGS_2020+REGS_2080;
  assign {FA_cout_3656,FA_out_3656}=REGS_1957+REGS_2021+REGS_2081;
  assign {FA_cout_3657,FA_out_3657}=REGS_1958+REGS_2022+REGS_2082;
  assign {FA_cout_3658,FA_out_3658}=REGS_1959+REGS_2023+REGS_2083;
  assign {FA_cout_3659,FA_out_3659}=REGS_1960+REGS_2024+REGS_2084;
  assign {FA_cout_3660,FA_out_3660}=REGS_1961+REGS_2025+REGS_2085;
  assign {FA_cout_3661,FA_out_3661}=REGS_1962+REGS_2026+REGS_2086;
  assign {FA_cout_3662,FA_out_3662}=REGS_1963+REGS_2027+REGS_2127;
  assign {FA_cout_3663,FA_out_3663}=REGS_2028+REGS_2029+REGS_2131;
  assign {FA_cout_3664,FA_out_3664}=REGS_2030+REGS_2031+REGS_2135;
  assign {FA_cout_3665,FA_out_3665}=REGS_2032+REGS_2033+REGS_2139;
  assign {FA_cout_3666,FA_out_3666}=REGS_2034+REGS_2035+REGS_2143;
  assign {FA_cout_3667,FA_out_3667}=REGS_2036+REGS_2037+REGS_2147;
  assign {FA_cout_3668,FA_out_3668}=REGS_2038+REGS_2087+REGS_2151;
  assign {FA_cout_3669,FA_out_3669}=REGS_2088+REGS_2128+REGS_2155;
  assign {FA_cout_3670,FA_out_3670}=REGS_2110+REGS_2262+REGS_2282;
  assign {FA_cout_3671,FA_out_3671}=REGS_2111+REGS_2263+REGS_2283;
  assign {FA_cout_3672,FA_out_3672}=REGS_2112+REGS_2264+REGS_2284;
  assign {FA_cout_3673,FA_out_3673}=REGS_2113+REGS_2265+REGS_2285;
  assign {FA_cout_3674,FA_out_3674}=REGS_2114+REGS_2266+REGS_2286;
  assign {FA_cout_3675,FA_out_3675}=REGS_2115+REGS_2267+REGS_2287;
  assign {FA_cout_3676,FA_out_3676}=REGS_2116+REGS_2268+REGS_2288;
  assign {FA_cout_3677,FA_out_3677}=REGS_2117+REGS_2269+REGS_2289;
  assign {FA_cout_3678,FA_out_3678}=REGS_2118+REGS_2270+REGS_2290;
  assign {FA_cout_3679,FA_out_3679}=REGS_2119+REGS_2271+REGS_2291;
  assign {FA_cout_3680,FA_out_3680}=REGS_2120+REGS_2272+REGS_2292;
  assign {FA_cout_3681,FA_out_3681}=REGS_2121+REGS_2273+REGS_2293;
  assign {FA_cout_3682,FA_out_3682}=REGS_2122+REGS_2274+REGS_2294;
  assign {FA_cout_3683,FA_out_3683}=REGS_2123+REGS_2275+REGS_2295;
  assign {FA_cout_3684,FA_out_3684}=REGS_2124+REGS_2276+REGS_2296;
  assign {FA_cout_3685,FA_out_3685}=REGS_2125+REGS_2277+REGS_2297;
  assign {FA_cout_3686,FA_out_3686}=REGS_2126+REGS_2278+REGS_2298;
  assign {FA_cout_3687,FA_out_3687}=REGS_2129+REGS_2132+REGS_2159;
  assign {FA_cout_3688,FA_out_3688}=REGS_2130+REGS_2299+REGS_2303;
  assign {FA_cout_3689,FA_out_3689}=REGS_2133+REGS_2136+REGS_2163;
  assign {FA_cout_3690,FA_out_3690}=REGS_2134+REGS_2304+REGS_2308;
  assign {FA_cout_3691,FA_out_3691}=REGS_2137+REGS_2140+REGS_2167;
  assign {FA_cout_3692,FA_out_3692}=REGS_2138+REGS_2309+REGS_2313;
  assign {FA_cout_3693,FA_out_3693}=REGS_2141+REGS_2144+REGS_2171;
  assign {FA_cout_3694,FA_out_3694}=REGS_2142+REGS_2314+REGS_2318;
  assign {FA_cout_3695,FA_out_3695}=REGS_2145+REGS_2148+REGS_2175;
  assign {FA_cout_3696,FA_out_3696}=REGS_2146+REGS_2319+REGS_2323;
  assign {FA_cout_3697,FA_out_3697}=REGS_2149+REGS_2152+REGS_2179;
  assign {FA_cout_3698,FA_out_3698}=REGS_2150+REGS_2324+REGS_2328;
  assign {FA_cout_3699,FA_out_3699}=REGS_2153+REGS_2156+REGS_2183;
  assign {FA_cout_3700,FA_out_3700}=REGS_2154+REGS_2329+REGS_2333;
  assign {FA_cout_3701,FA_out_3701}=REGS_2157+REGS_2160+REGS_2187;
  assign {FA_cout_3702,FA_out_3702}=REGS_2158+REGS_2334+REGS_2338;
  assign {FA_cout_3703,FA_out_3703}=REGS_2161+REGS_2164+REGS_2191;
  assign {FA_cout_3704,FA_out_3704}=REGS_2162+REGS_2339+REGS_2342;
  assign {FA_cout_3705,FA_out_3705}=REGS_2165+REGS_2168+REGS_2195;
  assign {FA_cout_3706,FA_out_3706}=REGS_2166+REGS_2343+REGS_2346;
  assign {FA_cout_3707,FA_out_3707}=REGS_2169+REGS_2172+REGS_2199;
  assign {FA_cout_3708,FA_out_3708}=REGS_2170+REGS_2347+REGS_2350;
  assign {FA_cout_3709,FA_out_3709}=REGS_2173+REGS_2176+REGS_2203;
  assign {FA_cout_3710,FA_out_3710}=REGS_2174+REGS_2351+REGS_2356;
  assign {FA_cout_3711,FA_out_3711}=REGS_2177+REGS_2180+REGS_2207;
  assign {FA_cout_3712,FA_out_3712}=REGS_2181+REGS_2184+REGS_2211;
  assign {FA_cout_3713,FA_out_3713}=REGS_2185+REGS_2188+REGS_2215;
  assign {FA_cout_3714,FA_out_3714}=REGS_2189+REGS_2192+REGS_2219;
  assign {FA_cout_3715,FA_out_3715}=REGS_2193+REGS_2196+REGS_2223;
  assign {FA_cout_3716,FA_out_3716}=REGS_2197+REGS_2200+REGS_2227;
  assign {FA_cout_3717,FA_out_3717}=REGS_2201+REGS_2204+REGS_2231;
  assign {FA_cout_3718,FA_out_3718}=REGS_2205+REGS_2208+REGS_2235;
  assign {FA_cout_3719,FA_out_3719}=REGS_2209+REGS_2212+REGS_2239;
  assign {FA_cout_3720,FA_out_3720}=REGS_2213+REGS_2216+REGS_2243;
  assign {FA_cout_3721,FA_out_3721}=REGS_2217+REGS_2220+REGS_2247;
  assign {FA_cout_3722,FA_out_3722}=REGS_2221+REGS_2224+REGS_2251;
  assign {FA_cout_3723,FA_out_3723}=REGS_2225+REGS_2228+REGS_2300;
  assign {FA_cout_3724,FA_out_3724}=REGS_2229+REGS_2232+REGS_2305;
  assign {FA_cout_3725,FA_out_3725}=REGS_2233+REGS_2236+REGS_2310;
  assign {FA_cout_3726,FA_out_3726}=REGS_2237+REGS_2240+REGS_2315;
  assign {FA_cout_3727,FA_out_3727}=REGS_2241+REGS_2244+REGS_2320;
  assign {FA_cout_3728,FA_out_3728}=REGS_2245+REGS_2248+REGS_2325;
  assign {FA_cout_3729,FA_out_3729}=REGS_2249+REGS_2252+REGS_2330;
  assign {FA_cout_3730,FA_out_3730}=REGS_2253+REGS_2280+REGS_2335;
  assign {FA_cout_3731,FA_out_3731}=FA_cout_3623+FA_out_3624+REGS_2089;
  assign {FA_cout_3732,FA_out_3732}=FA_cout_3624+FA_out_3625+REGS_2090;
  assign {FA_cout_3733,FA_out_3733}=FA_cout_3625+FA_out_3626+REGS_2091;
  assign {FA_cout_3734,FA_out_3734}=FA_cout_3626+FA_out_3627+REGS_2092;
  assign {FA_cout_3735,FA_out_3735}=FA_cout_3627+FA_out_3628+REGS_2093;
  assign {FA_cout_3736,FA_out_3736}=FA_cout_3628+FA_out_3629+REGS_2094;
  assign {FA_cout_3737,FA_out_3737}=FA_cout_3629+FA_out_3630+REGS_2095;
  assign {FA_cout_3738,FA_out_3738}=FA_cout_3630+FA_out_3631+REGS_2096;
  assign {FA_cout_3739,FA_out_3739}=FA_cout_3631+FA_out_3632+REGS_2097;
  assign {FA_cout_3740,FA_out_3740}=FA_cout_3632+FA_out_3633+REGS_2098;
  assign {FA_cout_3741,FA_out_3741}=FA_cout_3633+FA_out_3634+REGS_2099;
  assign {FA_cout_3742,FA_out_3742}=FA_cout_3634+FA_out_3635+REGS_2100;
  assign {FA_cout_3743,FA_out_3743}=FA_cout_3635+FA_out_3636+REGS_2101;
  assign {FA_cout_3744,FA_out_3744}=FA_cout_3636+FA_out_3637+HA_out_282;
  assign {FA_cout_3745,FA_out_3745}=FA_cout_3637+FA_out_3638+HA_cout_282;
  assign {FA_cout_3746,FA_out_3746}=FA_cout_3638+FA_out_3639+HA_cout_283;
  assign {FA_cout_3747,FA_out_3747}=FA_cout_3639+FA_out_3640+HA_cout_284;
  assign {FA_cout_3748,FA_out_3748}=FA_cout_3640+FA_out_3641+HA_cout_285;
  assign {FA_cout_3749,FA_out_3749}=FA_cout_3641+FA_out_3642+HA_cout_286;
  assign {FA_cout_3750,FA_out_3750}=FA_cout_3642+FA_out_3643+HA_cout_287;
  assign {FA_cout_3751,FA_out_3751}=FA_cout_3643+FA_out_3644+HA_cout_288;
  assign {FA_cout_3752,FA_out_3752}=FA_cout_3644+FA_out_3645+HA_cout_289;
  assign {FA_cout_3753,FA_out_3753}=FA_cout_3645+FA_out_3646+FA_cout_3670;
  assign {FA_cout_3754,FA_out_3754}=FA_cout_3646+FA_out_3647+FA_cout_3671;
  assign {FA_cout_3755,FA_out_3755}=FA_cout_3647+FA_out_3648+FA_cout_3672;
  assign {FA_cout_3756,FA_out_3756}=FA_cout_3648+FA_out_3649+FA_cout_3673;
  assign {FA_cout_3757,FA_out_3757}=FA_cout_3649+FA_out_3650+FA_cout_3674;
  assign {FA_cout_3758,FA_out_3758}=FA_cout_3650+FA_out_3651+FA_cout_3675;
  assign {FA_cout_3759,FA_out_3759}=FA_cout_3651+FA_out_3652+FA_cout_3676;
  assign {FA_cout_3760,FA_out_3760}=FA_cout_3652+FA_out_3653+FA_cout_3677;
  assign {FA_cout_3761,FA_out_3761}=FA_cout_3653+FA_out_3654+FA_cout_3678;
  assign {FA_cout_3762,FA_out_3762}=FA_cout_3654+FA_out_3655+FA_cout_3679;
  assign {FA_cout_3763,FA_out_3763}=FA_cout_3655+FA_out_3656+FA_cout_3680;
  assign {FA_cout_3764,FA_out_3764}=FA_cout_3656+FA_out_3657+FA_cout_3681;
  assign {FA_cout_3765,FA_out_3765}=FA_cout_3657+FA_out_3658+FA_cout_3682;
  assign {FA_cout_3766,FA_out_3766}=FA_cout_3658+FA_out_3659+FA_cout_3683;
  assign {FA_cout_3767,FA_out_3767}=FA_cout_3659+FA_out_3660+FA_cout_3684;
  assign {FA_cout_3768,FA_out_3768}=FA_cout_3660+FA_out_3661+FA_cout_3685;
  assign {FA_cout_3769,FA_out_3769}=FA_cout_3661+FA_out_3662+FA_cout_3686;
  assign {FA_cout_3770,FA_out_3770}=FA_cout_3662+FA_out_3663+FA_cout_3688;
  assign {FA_cout_3771,FA_out_3771}=FA_cout_3663+FA_out_3664+FA_cout_3690;
  assign {FA_cout_3772,FA_out_3772}=FA_cout_3664+FA_out_3665+FA_cout_3692;
  assign {FA_cout_3773,FA_out_3773}=FA_cout_3665+FA_out_3666+FA_cout_3694;
  assign {FA_cout_3774,FA_out_3774}=FA_cout_3666+FA_out_3667+FA_cout_3696;
  assign {FA_cout_3775,FA_out_3775}=FA_cout_3667+FA_out_3668+FA_cout_3698;
  assign {FA_cout_3776,FA_out_3776}=FA_cout_3668+FA_out_3669+FA_cout_3700;
  assign {FA_cout_3777,FA_out_3777}=FA_cout_3669+FA_out_3687+FA_cout_3702;
  assign {FA_cout_3778,FA_out_3778}=FA_cout_3687+FA_out_3689+FA_cout_3704;
  assign {FA_cout_3779,FA_out_3779}=FA_cout_3689+FA_out_3691+FA_cout_3706;
  assign {FA_cout_3780,FA_out_3780}=FA_cout_3691+FA_out_3693+FA_cout_3708;
  assign {FA_cout_3781,FA_out_3781}=FA_cout_3693+FA_out_3695+FA_cout_3710;
  assign {FA_cout_3782,FA_out_3782}=FA_cout_3695+FA_out_3697+HA_cout_290;
  assign {FA_cout_3783,FA_out_3783}=FA_cout_3697+FA_out_3699+HA_cout_291;
  assign {FA_cout_3784,FA_out_3784}=FA_cout_3699+FA_out_3701+HA_cout_292;
  assign {FA_cout_3785,FA_out_3785}=FA_cout_3701+FA_out_3703+HA_cout_293;
  assign {FA_cout_3786,FA_out_3786}=FA_cout_3703+FA_out_3705+HA_cout_294;
  assign {FA_cout_3787,FA_out_3787}=FA_cout_3705+FA_out_3707+HA_cout_295;
  assign {FA_cout_3788,FA_out_3788}=FA_cout_3707+FA_out_3709+REGS_2206;
  assign {FA_cout_3789,FA_out_3789}=FA_cout_3709+FA_out_3711+REGS_2210;
  assign {FA_cout_3790,FA_out_3790}=FA_cout_3711+FA_out_3712+REGS_2214;
  assign {FA_cout_3791,FA_out_3791}=FA_cout_3712+FA_out_3713+REGS_2218;
  assign {FA_cout_3792,FA_out_3792}=FA_cout_3713+FA_out_3714+REGS_2222;
  assign {FA_cout_3793,FA_out_3793}=FA_cout_3714+FA_out_3715+REGS_2226;
  assign {FA_cout_3794,FA_out_3794}=FA_cout_3715+FA_out_3716+REGS_2230;
  assign {FA_cout_3795,FA_out_3795}=FA_cout_3716+FA_out_3717+REGS_2234;
  assign {FA_cout_3796,FA_out_3796}=FA_cout_3717+FA_out_3718+REGS_2238;
  assign {FA_cout_3797,FA_out_3797}=FA_cout_3718+FA_out_3719+REGS_2242;
  assign {FA_cout_3798,FA_out_3798}=FA_cout_3719+FA_out_3720+REGS_2246;
  assign {FA_cout_3799,FA_out_3799}=FA_cout_3720+FA_out_3721+REGS_2250;
  assign {FA_cout_3800,FA_out_3800}=FA_cout_3721+FA_out_3722+REGS_2279;
  assign {FA_cout_3801,FA_out_3801}=FA_cout_3744+FA_out_3745+HA_out_283;
  assign {FA_cout_3802,FA_out_3802}=FA_cout_3745+FA_out_3746+HA_out_284;
  assign {FA_cout_3803,FA_out_3803}=FA_cout_3746+FA_out_3747+HA_out_285;
  assign {FA_cout_3804,FA_out_3804}=FA_cout_3747+FA_out_3748+HA_out_286;
  assign {FA_cout_3805,FA_out_3805}=FA_cout_3748+FA_out_3749+HA_out_287;
  assign {FA_cout_3806,FA_out_3806}=FA_cout_3749+FA_out_3750+HA_out_288;
  assign {FA_cout_3807,FA_out_3807}=FA_cout_3750+FA_out_3751+HA_out_289;
  assign {FA_cout_3808,FA_out_3808}=FA_cout_3751+FA_out_3752+FA_out_3670;
  assign {FA_cout_3809,FA_out_3809}=FA_cout_3752+FA_out_3753+FA_out_3671;
  assign {FA_cout_3810,FA_out_3810}=FA_cout_3753+FA_out_3754+FA_out_3672;
  assign {FA_cout_3811,FA_out_3811}=FA_cout_3754+FA_out_3755+FA_out_3673;
  assign {FA_cout_3812,FA_out_3812}=FA_cout_3755+FA_out_3756+FA_out_3674;
  assign {FA_cout_3813,FA_out_3813}=FA_cout_3756+FA_out_3757+FA_out_3675;
  assign {FA_cout_3814,FA_out_3814}=FA_cout_3757+FA_out_3758+FA_out_3676;
  assign {FA_cout_3815,FA_out_3815}=FA_cout_3758+FA_out_3759+FA_out_3677;
  assign {FA_cout_3816,FA_out_3816}=FA_cout_3759+FA_out_3760+FA_out_3678;
  assign {FA_cout_3817,FA_out_3817}=FA_cout_3760+FA_out_3761+FA_out_3679;
  assign {FA_cout_3818,FA_out_3818}=FA_cout_3761+FA_out_3762+FA_out_3680;
  assign {FA_cout_3819,FA_out_3819}=FA_cout_3762+FA_out_3763+FA_out_3681;
  assign {FA_cout_3820,FA_out_3820}=FA_cout_3763+FA_out_3764+FA_out_3682;
  assign {FA_cout_3821,FA_out_3821}=FA_cout_3764+FA_out_3765+HA_out_339;
  assign {FA_cout_3822,FA_out_3822}=FA_cout_3765+FA_out_3766+HA_cout_339;
  assign {FA_cout_3823,FA_out_3823}=FA_cout_3766+FA_out_3767+HA_cout_340;
  assign {FA_cout_3824,FA_out_3824}=FA_cout_3767+FA_out_3768+FA_out_3686;
  assign {FA_cout_3825,FA_out_3825}=FA_cout_3768+FA_out_3769+FA_out_3688;
  assign {FA_cout_3826,FA_out_3826}=FA_cout_3769+FA_out_3770+FA_out_3690;
  assign {FA_cout_3827,FA_out_3827}=FA_cout_3770+FA_out_3771+FA_out_3692;
  assign {FA_cout_3828,FA_out_3828}=FA_cout_3771+FA_out_3772+FA_out_3694;
  assign {FA_cout_3829,FA_out_3829}=FA_cout_3772+FA_out_3773+FA_out_3696;
  assign {FA_cout_3830,FA_out_3830}=FA_cout_3773+FA_out_3774+FA_out_3698;
  assign {FA_cout_3831,FA_out_3831}=FA_cout_3774+FA_out_3775+FA_out_3700;
  assign {FA_cout_3832,FA_out_3832}=FA_cout_3775+FA_out_3776+FA_out_3702;
  assign {FA_cout_3833,FA_out_3833}=FA_cout_3776+FA_out_3777+FA_out_3704;
  assign {FA_cout_3834,FA_out_3834}=FA_cout_3777+FA_out_3778+FA_out_3706;
  assign {FA_cout_3835,FA_out_3835}=FA_cout_3778+FA_out_3779+FA_out_3708;
  assign {FA_cout_3836,FA_out_3836}=FA_cout_3779+FA_out_3780+FA_out_3710;
  assign {FA_cout_3837,FA_out_3837}=FA_cout_3780+FA_out_3781+HA_out_290;
  assign {FA_cout_3838,FA_out_3838}=FA_cout_3781+FA_out_3782+HA_out_291;
  assign {FA_cout_3839,FA_out_3839}=FA_cout_3782+FA_out_3783+HA_out_292;
  assign {FA_cout_3840,FA_out_3840}=FA_cout_3783+FA_out_3784+HA_out_293;
  assign {FA_cout_3841,FA_out_3841}=FA_cout_3784+FA_out_3785+HA_out_294;
  assign {FA_cout_3842,FA_out_3842}=FA_cout_3785+FA_out_3786+HA_out_295;
  assign {FA_cout_3843,FA_out_3843}=FA_cout_3786+FA_out_3787+REGS_2202;
  assign {FA_cout_3844,FA_out_3844}=FA_cout_3821+FA_out_3822+HA_out_340;
  assign {FA_cout_3845,FA_out_3845}=FA_cout_3822+FA_out_3823+FA_out_3685;
  assign {HA_cout_0,HA_out_0}=inp_0[1]+inp_1[0];
  assign {HA_cout_1,HA_out_1}=inp_3[1]+inp_4[0];
  assign {HA_cout_2,HA_out_2}=inp_6[1]+inp_7[0];
  assign {HA_cout_3,HA_out_3}=inp_9[1]+inp_10[0];
  assign {HA_cout_4,HA_out_4}=inp_12[1]+inp_13[0];
  assign {HA_cout_5,HA_out_5}=inp_15[1]+inp_16[0];
  assign {HA_cout_6,HA_out_6}=inp_18[1]+inp_19[0];
  assign {HA_cout_7,HA_out_7}=inp_21[1]+inp_22[0];
  assign {HA_cout_8,HA_out_8}=inp_24[1]+inp_25[0];
  assign {HA_cout_9,HA_out_9}=inp_27[1]+inp_28[0];
  assign {HA_cout_10,HA_out_10}=inp_30[1]+inp_31[0];
  assign {HA_cout_11,HA_out_11}=inp_33[1]+inp_34[0];
  assign {HA_cout_12,HA_out_12}=inp_36[1]+inp_37[0];
  assign {HA_cout_13,HA_out_13}=inp_39[1]+inp_40[0];
  assign {HA_cout_14,HA_out_14}=inp_42[1]+inp_43[0];
  assign {HA_cout_15,HA_out_15}=inp_45[1]+inp_46[0];
  assign {HA_cout_16,HA_out_16}=inp_48[1]+inp_49[0];
  assign {HA_cout_17,HA_out_17}=inp_51[1]+inp_52[0];
  assign {HA_cout_18,HA_out_18}=inp_54[1]+inp_55[0];
  assign {HA_cout_19,HA_out_19}=inp_57[1]+inp_58[0];
  assign {HA_cout_20,HA_out_20}=inp_60[1]+inp_61[0];
  assign {HA_cout_21,HA_out_21}=inp_62[3]+inp_63[2];
  assign {HA_cout_22,HA_out_22}=inp_62[6]+inp_63[5];
  assign {HA_cout_23,HA_out_23}=inp_62[9]+inp_63[8];
  assign {HA_cout_24,HA_out_24}=inp_62[12]+inp_63[11];
  assign {HA_cout_25,HA_out_25}=inp_62[15]+inp_63[14];
  assign {HA_cout_26,HA_out_26}=inp_62[18]+inp_63[17];
  assign {HA_cout_27,HA_out_27}=inp_62[21]+inp_63[20];
  assign {HA_cout_28,HA_out_28}=inp_62[24]+inp_63[23];
  assign {HA_cout_29,HA_out_29}=inp_62[27]+inp_63[26];
  assign {HA_cout_30,HA_out_30}=inp_62[30]+inp_63[29];
  assign {HA_cout_31,HA_out_31}=inp_62[33]+inp_63[32];
  assign {HA_cout_32,HA_out_32}=inp_62[36]+inp_63[35];
  assign {HA_cout_33,HA_out_33}=inp_62[39]+inp_63[38];
  assign {HA_cout_34,HA_out_34}=inp_62[42]+inp_63[41];
  assign {HA_cout_35,HA_out_35}=inp_62[45]+inp_63[44];
  assign {HA_cout_36,HA_out_36}=inp_62[48]+inp_63[47];
  assign {HA_cout_37,HA_out_37}=inp_62[51]+inp_63[50];
  assign {HA_cout_38,HA_out_38}=inp_62[54]+inp_63[53];
  assign {HA_cout_39,HA_out_39}=inp_62[57]+inp_63[56];
  assign {HA_cout_40,HA_out_40}=inp_62[60]+inp_63[59];
  assign {HA_cout_41,HA_out_41}=inp_62[63]+inp_63[62];
  assign {HA_cout_42,HA_out_42}=HA_cout_0+FA_out_0;
  assign {HA_cout_43,HA_out_43}=FA_out_65+inp_6[0];
  assign {HA_cout_44,HA_out_44}=FA_out_66+HA_out_2;
  assign {HA_cout_45,HA_out_45}=HA_cout_3+FA_out_192;
  assign {HA_cout_46,HA_out_46}=FA_out_257+inp_15[0];
  assign {HA_cout_47,HA_out_47}=FA_out_258+HA_out_5;
  assign {HA_cout_48,HA_out_48}=HA_cout_6+FA_out_384;
  assign {HA_cout_49,HA_out_49}=FA_out_449+inp_24[0];
  assign {HA_cout_50,HA_out_50}=FA_out_450+HA_out_8;
  assign {HA_cout_51,HA_out_51}=HA_cout_9+FA_out_576;
  assign {HA_cout_52,HA_out_52}=FA_out_640+sm_sig;
  assign {HA_cout_53,HA_out_53}=FA_out_641+inp_33[0];
  assign {HA_cout_54,HA_out_54}=FA_out_642+HA_out_11;
  assign {HA_cout_55,HA_out_55}=HA_cout_12+FA_out_768;
  assign {HA_cout_56,HA_out_56}=FA_out_833+inp_42[0];
  assign {HA_cout_57,HA_out_57}=FA_out_834+HA_out_14;
  assign {HA_cout_58,HA_out_58}=HA_cout_15+FA_out_960;
  assign {HA_cout_59,HA_out_59}=FA_out_1025+inp_51[0];
  assign {HA_cout_60,HA_out_60}=FA_out_1026+HA_out_17;
  assign {HA_cout_61,HA_out_61}=HA_cout_18+FA_out_1152;
  assign {HA_cout_62,HA_out_62}=FA_out_1217+inp_60[0];
  assign {HA_cout_63,HA_out_63}=FA_out_1218+HA_out_20;
  assign {HA_cout_64,HA_out_64}=FA_cout_1284+FA_out_1304;
  assign {HA_cout_65,HA_out_65}=FA_cout_1287+FA_out_1307;
  assign {HA_cout_66,HA_out_66}=FA_cout_1290+FA_out_1310;
  assign {HA_cout_67,HA_out_67}=FA_cout_1293+FA_out_1313;
  assign {HA_cout_68,HA_out_68}=FA_cout_1296+FA_out_1316;
  assign {HA_cout_69,HA_out_69}=FA_cout_1299+FA_out_1319;
  assign {HA_cout_70,HA_out_70}=FA_cout_1302+FA_out_1322;
  assign {HA_cout_71,HA_out_71}=FA_cout_1304+HA_out_23;
  assign {HA_cout_72,HA_out_72}=FA_cout_1307+HA_out_26;
  assign {HA_cout_73,HA_out_73}=FA_cout_1310+HA_out_29;
  assign {HA_cout_74,HA_out_74}=FA_cout_1313+HA_out_32;
  assign {HA_cout_75,HA_out_75}=FA_cout_1316+HA_out_35;
  assign {HA_cout_76,HA_out_76}=FA_cout_1319+HA_out_38;
  assign {HA_cout_77,HA_out_77}=FA_cout_1322+HA_out_41;
  assign {HA_cout_78,HA_out_78}=HA_cout_23+inp_63[9];
  assign {HA_cout_79,HA_out_79}=HA_cout_26+inp_63[18];
  assign {HA_cout_80,HA_out_80}=HA_cout_29+inp_63[27];
  assign {HA_cout_81,HA_out_81}=HA_cout_32+inp_63[36];
  assign {HA_cout_82,HA_out_82}=HA_cout_35+inp_63[45];
  assign {HA_cout_83,HA_out_83}=HA_cout_38+inp_63[54];
  assign {HA_cout_84,HA_out_84}=HA_cout_41+inp_63[63];
  assign {HA_cout_85,HA_out_85}=REGS_3+REGS_67;
  assign {HA_cout_86,HA_out_86}=REGS_4+REGS_68;
  assign {HA_cout_87,HA_out_87}=REGS_199+REGS_271;
  assign {HA_cout_88,HA_out_88}=REGS_200+REGS_272;
  assign {HA_cout_89,HA_out_89}=REGS_201+REGS_273;
  assign {HA_cout_90,HA_out_90}=REGS_405+REGS_461;
  assign {HA_cout_91,HA_out_91}=REGS_406+REGS_462;
  assign {HA_cout_92,HA_out_92}=REGS_601+REGS_672;
  assign {HA_cout_93,HA_out_93}=REGS_602+REGS_673;
  assign {HA_cout_94,HA_out_94}=REGS_816+REGS_865;
  assign {HA_cout_95,HA_out_95}=REGS_817+REGS_866;
  assign {HA_cout_96,HA_out_96}=REGS_992+REGS_1085;
  assign {HA_cout_97,HA_out_97}=REGS_993+REGS_1086;
  assign {HA_cout_98,HA_out_98}=REGS_994+REGS_1087;
  assign {HA_cout_99,HA_out_99}=REGS_1213+REGS_1254;
  assign {HA_cout_100,HA_out_100}=REGS_1214+REGS_1255;
  assign {HA_cout_101,HA_out_101}=REGS_1400+REGS_1480;
  assign {HA_cout_102,HA_out_102}=REGS_1401+REGS_1481;
  assign {HA_cout_103,HA_out_103}=REGS_1630+REGS_1664;
  assign {HA_cout_104,HA_out_104}=REGS_1631+REGS_1665;
  assign {HA_cout_105,HA_out_105}=REGS_1760+REGS_1866;
  assign {HA_cout_106,HA_out_106}=REGS_1763+REGS_1794;
  assign {HA_cout_107,HA_out_107}=REGS_1766+REGS_1871;
  assign {HA_cout_108,HA_out_108}=REGS_1772+REGS_1875;
  assign {HA_cout_109,HA_out_109}=REGS_1775+REGS_1806;
  assign {HA_cout_110,HA_out_110}=REGS_1778+REGS_1880;
  assign {HA_cout_111,HA_out_111}=REGS_1784+REGS_1884;
  assign {HA_cout_112,HA_out_112}=REGS_1785+REGS_1885;
  assign {HA_cout_113,HA_out_113}=REGS_1789+REGS_1816;
  assign {HA_cout_114,HA_out_114}=REGS_1792+REGS_1887;
  assign {HA_cout_115,HA_out_115}=REGS_1795+REGS_1822;
  assign {HA_cout_116,HA_out_116}=REGS_1801+REGS_1828;
  assign {HA_cout_117,HA_out_117}=REGS_1804+REGS_1890;
  assign {HA_cout_118,HA_out_118}=REGS_1807+REGS_1834;
  assign {HA_cout_119,HA_out_119}=REGS_1813+REGS_1840;
  assign {HA_cout_120,HA_out_120}=REGS_1817+REGS_1843;
  assign {HA_cout_121,HA_out_121}=REGS_1823+REGS_1848;
  assign {HA_cout_122,HA_out_122}=REGS_1829+REGS_1852;
  assign {HA_cout_123,HA_out_123}=REGS_1835+REGS_1857;
  assign {HA_cout_124,HA_out_124}=REGS_1841+REGS_1861;
  assign {HA_cout_125,HA_out_125}=REGS_1844+REGS_1864;
  assign {HA_cout_126,HA_out_126}=REGS_1853+REGS_1873;
  assign {HA_cout_127,HA_out_127}=REGS_1862+REGS_1882;
  assign {HA_cout_128,HA_out_128}=HA_cout_85+HA_out_86;
  assign {HA_cout_129,HA_out_129}=HA_cout_86+FA_out_2205;
  assign {HA_cout_130,HA_out_130}=FA_cout_2205+FA_out_2206;
  assign {HA_cout_131,HA_out_131}=FA_out_2272+REGS_403;
  assign {HA_cout_132,HA_out_132}=FA_out_2273+REGS_404;
  assign {HA_cout_133,HA_out_133}=FA_out_2274+HA_out_90;
  assign {HA_cout_134,HA_out_134}=HA_cout_92+HA_out_93;
  assign {HA_cout_135,HA_out_135}=HA_cout_93+FA_out_2404;
  assign {HA_cout_136,HA_out_136}=FA_cout_2404+FA_out_2405;
  assign {HA_cout_137,HA_out_137}=FA_out_2477+REGS_989;
  assign {HA_cout_138,HA_out_138}=FA_out_2478+REGS_990;
  assign {HA_cout_139,HA_out_139}=FA_out_2479+REGS_991;
  assign {HA_cout_140,HA_out_140}=FA_out_2480+HA_out_96;
  assign {HA_cout_141,HA_out_141}=HA_cout_99+HA_out_100;
  assign {HA_cout_142,HA_out_142}=HA_cout_100+FA_out_2608;
  assign {HA_cout_143,HA_out_143}=FA_cout_2608+FA_out_2609;
  assign {HA_cout_144,HA_out_144}=FA_cout_2609+FA_out_2610;
  assign {HA_cout_145,HA_out_145}=FA_out_2672+REGS_1627;
  assign {HA_cout_146,HA_out_146}=FA_out_2673+REGS_1628;
  assign {HA_cout_147,HA_out_147}=FA_out_2674+REGS_1629;
  assign {HA_cout_148,HA_out_148}=FA_out_2675+HA_out_103;
  assign {HA_cout_149,HA_out_149}=FA_cout_2759+FA_out_2767;
  assign {HA_cout_150,HA_out_150}=FA_out_2761+REGS_1891;
  assign {HA_cout_151,HA_out_151}=FA_out_2766+REGS_1826;
  assign {HA_cout_152,HA_out_152}=FA_cout_2767+FA_out_2776;
  assign {HA_cout_153,HA_out_153}=FA_cout_2773+FA_out_2782;
  assign {HA_cout_154,HA_out_154}=FA_out_2775+REGS_1851;
  assign {HA_cout_155,HA_out_155}=FA_cout_2776+FA_out_2785;
  assign {HA_cout_156,HA_out_156}=FA_cout_2779+FA_out_2788;
  assign {HA_cout_157,HA_out_157}=FA_cout_2782+HA_out_106;
  assign {HA_cout_158,HA_out_158}=FA_cout_2785+HA_out_108;
  assign {HA_cout_159,HA_out_159}=FA_cout_2788+FA_out_2791;
  assign {HA_cout_160,HA_out_160}=HA_cout_106+HA_out_115;
  assign {HA_cout_161,HA_out_161}=HA_cout_108+HA_out_117;
  assign {HA_cout_162,HA_out_162}=FA_cout_2791+HA_out_119;
  assign {HA_cout_163,HA_out_163}=HA_cout_111+HA_out_112;
  assign {HA_cout_164,HA_out_164}=HA_cout_112+REGS_1786;
  assign {HA_cout_165,HA_out_165}=HA_cout_115+HA_out_121;
  assign {HA_cout_166,HA_out_166}=HA_cout_117+REGS_1832;
  assign {HA_cout_167,HA_out_167}=HA_cout_119+HA_out_124;
  assign {HA_cout_168,HA_out_168}=HA_cout_121+REGS_1869;
  assign {HA_cout_169,HA_out_169}=HA_cout_124+HA_out_127;
  assign {HA_cout_170,HA_out_170}=HA_cout_127+REGS_1883;
  assign {HA_cout_171,HA_out_171}=HA_cout_128+HA_out_129;
  assign {HA_cout_172,HA_out_172}=HA_cout_129+HA_out_130;
  assign {HA_cout_173,HA_out_173}=HA_cout_130+FA_out_2792;
  assign {HA_cout_174,HA_out_174}=FA_cout_2792+FA_out_2793;
  assign {HA_cout_175,HA_out_175}=FA_cout_2793+FA_out_2794;
  assign {HA_cout_176,HA_out_176}=FA_out_2861+REGS_599;
  assign {HA_cout_177,HA_out_177}=FA_out_2862+REGS_600;
  assign {HA_cout_178,HA_out_178}=FA_out_2863+HA_out_92;
  assign {HA_cout_179,HA_out_179}=FA_out_2864+HA_out_134;
  assign {HA_cout_180,HA_out_180}=HA_cout_137+HA_out_138;
  assign {HA_cout_181,HA_out_181}=HA_cout_138+HA_out_139;
  assign {HA_cout_182,HA_out_182}=HA_cout_139+HA_out_140;
  assign {HA_cout_183,HA_out_183}=HA_cout_140+FA_out_2998;
  assign {HA_cout_184,HA_out_184}=FA_cout_2998+FA_out_2999;
  assign {HA_cout_185,HA_out_185}=FA_cout_2999+FA_out_3000;
  assign {HA_cout_186,HA_out_186}=FA_cout_3000+FA_out_3001;
  assign {HA_cout_187,HA_out_187}=FA_out_3078+HA_out_102;
  assign {HA_cout_188,HA_out_188}=FA_out_3079+FA_out_2670;
  assign {HA_cout_189,HA_out_189}=FA_out_3080+FA_out_2671;
  assign {HA_cout_190,HA_out_190}=FA_out_3081+HA_out_145;
  assign {HA_cout_191,HA_out_191}=FA_out_3146+REGS_1876;
  assign {HA_cout_192,HA_out_192}=FA_out_3149+FA_out_2772;
  assign {HA_cout_193,HA_out_193}=FA_cout_3150+FA_out_3156;
  assign {HA_cout_194,HA_out_194}=FA_out_3155+FA_out_2781;
  assign {HA_cout_195,HA_out_195}=FA_cout_3156+FA_out_3162;
  assign {HA_cout_196,HA_out_196}=FA_out_3161+HA_out_105;
  assign {HA_cout_197,HA_out_197}=FA_cout_3162+FA_out_3168;
  assign {HA_cout_198,HA_out_198}=FA_out_3167+HA_out_114;
  assign {HA_cout_199,HA_out_199}=FA_cout_3168+FA_out_3174;
  assign {HA_cout_200,HA_out_200}=FA_out_3173+REGS_1820;
  assign {HA_cout_201,HA_out_201}=FA_cout_3174+FA_out_3180;
  assign {HA_cout_202,HA_out_202}=FA_cout_3177+FA_out_3181;
  assign {HA_cout_203,HA_out_203}=FA_cout_3180+HA_out_151;
  assign {HA_cout_204,HA_out_204}=FA_cout_3181+FA_out_3183;
  assign {HA_cout_205,HA_out_205}=HA_cout_151+HA_out_154;
  assign {HA_cout_206,HA_out_206}=FA_cout_3183+HA_out_156;
  assign {HA_cout_207,HA_out_207}=HA_cout_154+FA_out_2784;
  assign {HA_cout_208,HA_out_208}=HA_cout_156+HA_out_159;
  assign {HA_cout_209,HA_out_209}=HA_cout_159+HA_out_162;
  assign {HA_cout_210,HA_out_210}=HA_cout_162+HA_out_167;
  assign {HA_cout_211,HA_out_211}=HA_cout_163+HA_out_164;
  assign {HA_cout_212,HA_out_212}=HA_cout_164+REGS_1814;
  assign {HA_cout_213,HA_out_213}=HA_cout_167+HA_out_169;
  assign {HA_cout_214,HA_out_214}=HA_cout_169+HA_out_170;
  assign {HA_cout_215,HA_out_215}=HA_cout_171+HA_out_172;
  assign {HA_cout_216,HA_out_216}=HA_cout_172+HA_out_173;
  assign {HA_cout_217,HA_out_217}=HA_cout_173+HA_out_174;
  assign {HA_cout_218,HA_out_218}=HA_cout_174+HA_out_175;
  assign {HA_cout_219,HA_out_219}=HA_cout_175+FA_out_3184;
  assign {HA_cout_220,HA_out_220}=FA_cout_3184+FA_out_3185;
  assign {HA_cout_221,HA_out_221}=FA_cout_3185+FA_out_3186;
  assign {HA_cout_222,HA_out_222}=FA_cout_3186+FA_out_3187;
  assign {HA_cout_223,HA_out_223}=FA_cout_3187+FA_out_3188;
  assign {HA_cout_224,HA_out_224}=FA_out_3254+HA_out_95;
  assign {HA_cout_225,HA_out_225}=FA_out_3255+FA_out_2476;
  assign {HA_cout_226,HA_out_226}=FA_out_3256+HA_out_137;
  assign {HA_cout_227,HA_out_227}=FA_out_3257+HA_out_180;
  assign {HA_cout_228,HA_out_228}=FA_out_3386+HA_out_116;
  assign {HA_cout_229,HA_out_229}=FA_out_3389+HA_out_122;
  assign {HA_cout_230,HA_out_230}=FA_out_3392+HA_out_126;
  assign {HA_cout_231,HA_out_231}=FA_out_3395+REGS_1874;
  assign {HA_cout_232,HA_out_232}=HA_cout_187+HA_out_188;
  assign {HA_cout_233,HA_out_233}=HA_cout_188+HA_out_189;
  assign {HA_cout_234,HA_out_234}=HA_cout_189+HA_out_190;
  assign {HA_cout_235,HA_out_235}=HA_cout_190+FA_out_3397;
  assign {HA_cout_236,HA_out_236}=FA_cout_3397+FA_out_3398;
  assign {HA_cout_237,HA_out_237}=FA_cout_3398+FA_out_3399;
  assign {HA_cout_238,HA_out_238}=FA_cout_3399+FA_out_3400;
  assign {HA_cout_239,HA_out_239}=FA_cout_3400+FA_out_3401;
  assign {HA_cout_240,HA_out_240}=FA_cout_3401+FA_out_3402;
  assign {HA_cout_241,HA_out_241}=FA_cout_3409+FA_out_3413;
  assign {HA_cout_242,HA_out_242}=FA_cout_3413+FA_out_3417;
  assign {HA_cout_243,HA_out_243}=FA_cout_3417+FA_out_3421;
  assign {HA_cout_244,HA_out_244}=FA_cout_3421+FA_out_3425;
  assign {HA_cout_245,HA_out_245}=FA_cout_3425+FA_out_3429;
  assign {HA_cout_246,HA_out_246}=FA_cout_3429+FA_out_3433;
  assign {HA_cout_247,HA_out_247}=FA_cout_3433+FA_out_3437;
  assign {HA_cout_248,HA_out_248}=FA_cout_3437+HA_out_192;
  assign {HA_cout_249,HA_out_249}=FA_cout_3439+FA_out_3440;
  assign {HA_cout_250,HA_out_250}=HA_cout_192+HA_out_194;
  assign {HA_cout_251,HA_out_251}=FA_cout_3440+FA_out_3441;
  assign {HA_cout_252,HA_out_252}=HA_cout_194+HA_out_196;
  assign {HA_cout_253,HA_out_253}=FA_cout_3441+FA_out_3442;
  assign {HA_cout_254,HA_out_254}=HA_cout_196+HA_out_198;
  assign {HA_cout_255,HA_out_255}=FA_cout_3442+FA_out_3443;
  assign {HA_cout_256,HA_out_256}=HA_cout_198+HA_out_200;
  assign {HA_cout_257,HA_out_257}=FA_cout_3443+HA_out_202;
  assign {HA_cout_258,HA_out_258}=HA_cout_200+FA_out_3179;
  assign {HA_cout_259,HA_out_259}=HA_cout_202+HA_out_204;
  assign {HA_cout_260,HA_out_260}=HA_cout_204+HA_out_206;
  assign {HA_cout_261,HA_out_261}=HA_cout_206+HA_out_208;
  assign {HA_cout_262,HA_out_262}=HA_cout_208+HA_out_209;
  assign {HA_cout_263,HA_out_263}=HA_cout_209+HA_out_210;
  assign {HA_cout_264,HA_out_264}=HA_cout_210+HA_out_213;
  assign {HA_cout_265,HA_out_265}=HA_cout_213+HA_out_214;
  assign {HA_cout_266,HA_out_266}=HA_cout_214+HA_cout_170;
  assign {HA_cout_267,HA_out_267}=REGS_1900+REGS_1964;
  assign {HA_cout_268,HA_out_268}=REGS_1901+REGS_1965;
  assign {HA_cout_269,HA_out_269}=REGS_1902+REGS_1966;
  assign {HA_cout_270,HA_out_270}=REGS_1903+REGS_1967;
  assign {HA_cout_271,HA_out_271}=REGS_1904+REGS_1968;
  assign {HA_cout_272,HA_out_272}=REGS_1905+REGS_1969;
  assign {HA_cout_273,HA_out_273}=REGS_1906+REGS_1970;
  assign {HA_cout_274,HA_out_274}=REGS_1907+REGS_1971;
  assign {HA_cout_275,HA_out_275}=REGS_1908+REGS_1972;
  assign {HA_cout_276,HA_out_276}=REGS_1909+REGS_1973;
  assign {HA_cout_277,HA_out_277}=REGS_1910+REGS_1974;
  assign {HA_cout_278,HA_out_278}=REGS_1911+REGS_1975;
  assign {HA_cout_279,HA_out_279}=REGS_1912+REGS_1976;
  assign {HA_cout_280,HA_out_280}=REGS_1913+REGS_1977;
  assign {HA_cout_281,HA_out_281}=REGS_1914+REGS_1978;
  assign {HA_cout_282,HA_out_282}=REGS_2102+REGS_2254;
  assign {HA_cout_283,HA_out_283}=REGS_2103+REGS_2255;
  assign {HA_cout_284,HA_out_284}=REGS_2104+REGS_2256;
  assign {HA_cout_285,HA_out_285}=REGS_2105+REGS_2257;
  assign {HA_cout_286,HA_out_286}=REGS_2106+REGS_2258;
  assign {HA_cout_287,HA_out_287}=REGS_2107+REGS_2259;
  assign {HA_cout_288,HA_out_288}=REGS_2108+REGS_2260;
  assign {HA_cout_289,HA_out_289}=REGS_2109+REGS_2261;
  assign {HA_cout_290,HA_out_290}=REGS_2178+REGS_2359;
  assign {HA_cout_291,HA_out_291}=REGS_2182+REGS_2362;
  assign {HA_cout_292,HA_out_292}=REGS_2186+REGS_2365;
  assign {HA_cout_293,HA_out_293}=REGS_2190+REGS_2368;
  assign {HA_cout_294,HA_out_294}=REGS_2194+REGS_2372;
  assign {HA_cout_295,HA_out_295}=REGS_2198+REGS_2376;
  assign {HA_cout_296,HA_out_296}=REGS_2281+REGS_2301;
  assign {HA_cout_297,HA_out_297}=REGS_2302+REGS_2306;
  assign {HA_cout_298,HA_out_298}=REGS_2307+REGS_2311;
  assign {HA_cout_299,HA_out_299}=REGS_2312+REGS_2316;
  assign {HA_cout_300,HA_out_300}=REGS_2317+REGS_2321;
  assign {HA_cout_301,HA_out_301}=REGS_2322+REGS_2326;
  assign {HA_cout_302,HA_out_302}=REGS_2327+REGS_2331;
  assign {HA_cout_303,HA_out_303}=REGS_2332+REGS_2336;
  assign {HA_cout_304,HA_out_304}=REGS_2337+REGS_2340;
  assign {HA_cout_305,HA_out_305}=REGS_2341+REGS_2344;
  assign {HA_cout_306,HA_out_306}=REGS_2345+REGS_2348;
  assign {HA_cout_307,HA_out_307}=REGS_2349+REGS_2352;
  assign {HA_cout_308,HA_out_308}=REGS_2353+REGS_2354;
  assign {HA_cout_309,HA_out_309}=REGS_2355+REGS_2357;
  assign {HA_cout_310,HA_out_310}=REGS_2358+REGS_2360;
  assign {HA_cout_311,HA_out_311}=REGS_2361+REGS_2363;
  assign {HA_cout_312,HA_out_312}=REGS_2364+REGS_2366;
  assign {HA_cout_313,HA_out_313}=REGS_2367+REGS_2369;
  assign {HA_cout_314,HA_out_314}=REGS_2370+REGS_2373;
  assign {HA_cout_315,HA_out_315}=HA_cout_267+HA_out_268;
  assign {HA_cout_316,HA_out_316}=HA_cout_268+HA_out_269;
  assign {HA_cout_317,HA_out_317}=HA_cout_269+HA_out_270;
  assign {HA_cout_318,HA_out_318}=HA_cout_270+HA_out_271;
  assign {HA_cout_319,HA_out_319}=HA_cout_271+HA_out_272;
  assign {HA_cout_320,HA_out_320}=HA_cout_272+HA_out_273;
  assign {HA_cout_321,HA_out_321}=HA_cout_273+HA_out_274;
  assign {HA_cout_322,HA_out_322}=HA_cout_274+HA_out_275;
  assign {HA_cout_323,HA_out_323}=HA_cout_275+HA_out_276;
  assign {HA_cout_324,HA_out_324}=HA_cout_276+HA_out_277;
  assign {HA_cout_325,HA_out_325}=HA_cout_277+HA_out_278;
  assign {HA_cout_326,HA_out_326}=HA_cout_278+HA_out_279;
  assign {HA_cout_327,HA_out_327}=HA_cout_279+HA_out_280;
  assign {HA_cout_328,HA_out_328}=HA_cout_280+HA_out_281;
  assign {HA_cout_329,HA_out_329}=HA_cout_281+FA_out_3614;
  assign {HA_cout_330,HA_out_330}=FA_cout_3614+FA_out_3615;
  assign {HA_cout_331,HA_out_331}=FA_cout_3615+FA_out_3616;
  assign {HA_cout_332,HA_out_332}=FA_cout_3616+FA_out_3617;
  assign {HA_cout_333,HA_out_333}=FA_cout_3617+FA_out_3618;
  assign {HA_cout_334,HA_out_334}=FA_cout_3618+FA_out_3619;
  assign {HA_cout_335,HA_out_335}=FA_cout_3619+FA_out_3620;
  assign {HA_cout_336,HA_out_336}=FA_cout_3620+FA_out_3621;
  assign {HA_cout_337,HA_out_337}=FA_cout_3621+FA_out_3622;
  assign {HA_cout_338,HA_out_338}=FA_cout_3622+FA_out_3623;
  assign {HA_cout_339,HA_out_339}=FA_out_3683+REGS_2371;
  assign {HA_cout_340,HA_out_340}=FA_out_3684+REGS_2375;
  assign {HA_cout_341,HA_out_341}=FA_cout_3722+FA_out_3723;
  assign {HA_cout_342,HA_out_342}=FA_cout_3723+FA_out_3724;
  assign {HA_cout_343,HA_out_343}=FA_cout_3724+FA_out_3725;
  assign {HA_cout_344,HA_out_344}=FA_cout_3725+FA_out_3726;
  assign {HA_cout_345,HA_out_345}=FA_cout_3726+FA_out_3727;
  assign {HA_cout_346,HA_out_346}=FA_cout_3727+FA_out_3728;
  assign {HA_cout_347,HA_out_347}=FA_cout_3728+FA_out_3729;
  assign {HA_cout_348,HA_out_348}=FA_cout_3729+FA_out_3730;
  assign {HA_cout_349,HA_out_349}=FA_cout_3730+HA_out_296;
  assign {HA_cout_350,HA_out_350}=HA_cout_296+HA_out_297;
  assign {HA_cout_351,HA_out_351}=HA_cout_297+HA_out_298;
  assign {HA_cout_352,HA_out_352}=HA_cout_298+HA_out_299;
  assign {HA_cout_353,HA_out_353}=HA_cout_299+HA_out_300;
  assign {HA_cout_354,HA_out_354}=HA_cout_300+HA_out_301;
  assign {HA_cout_355,HA_out_355}=HA_cout_301+HA_out_302;
  assign {HA_cout_356,HA_out_356}=HA_cout_302+HA_out_303;
  assign {HA_cout_357,HA_out_357}=HA_cout_303+HA_out_304;
  assign {HA_cout_358,HA_out_358}=HA_cout_304+HA_out_305;
  assign {HA_cout_359,HA_out_359}=HA_cout_305+HA_out_306;
  assign {HA_cout_360,HA_out_360}=HA_cout_306+HA_out_307;
  assign {HA_cout_361,HA_out_361}=HA_cout_307+HA_out_308;
  assign {HA_cout_362,HA_out_362}=HA_cout_308+HA_out_309;
  assign {HA_cout_363,HA_out_363}=HA_cout_309+HA_out_310;
  assign {HA_cout_364,HA_out_364}=HA_cout_310+HA_out_311;
  assign {HA_cout_365,HA_out_365}=HA_cout_311+HA_out_312;
  assign {HA_cout_366,HA_out_366}=HA_cout_312+HA_out_313;
  assign {HA_cout_367,HA_out_367}=HA_cout_313+HA_out_314;
  assign {HA_cout_368,HA_out_368}=HA_cout_314+REGS_2374;
  assign {HA_cout_369,HA_out_369}=HA_cout_315+HA_out_316;
  assign {HA_cout_370,HA_out_370}=HA_cout_316+HA_out_317;
  assign {HA_cout_371,HA_out_371}=HA_cout_317+HA_out_318;
  assign {HA_cout_372,HA_out_372}=HA_cout_318+HA_out_319;
  assign {HA_cout_373,HA_out_373}=HA_cout_319+HA_out_320;
  assign {HA_cout_374,HA_out_374}=HA_cout_320+HA_out_321;
  assign {HA_cout_375,HA_out_375}=HA_cout_321+HA_out_322;
  assign {HA_cout_376,HA_out_376}=HA_cout_322+HA_out_323;
  assign {HA_cout_377,HA_out_377}=HA_cout_323+HA_out_324;
  assign {HA_cout_378,HA_out_378}=HA_cout_324+HA_out_325;
  assign {HA_cout_379,HA_out_379}=HA_cout_325+HA_out_326;
  assign {HA_cout_380,HA_out_380}=HA_cout_326+HA_out_327;
  assign {HA_cout_381,HA_out_381}=HA_cout_327+HA_out_328;
  assign {HA_cout_382,HA_out_382}=HA_cout_328+HA_out_329;
  assign {HA_cout_383,HA_out_383}=HA_cout_329+HA_out_330;
  assign {HA_cout_384,HA_out_384}=HA_cout_330+HA_out_331;
  assign {HA_cout_385,HA_out_385}=HA_cout_331+HA_out_332;
  assign {HA_cout_386,HA_out_386}=HA_cout_332+HA_out_333;
  assign {HA_cout_387,HA_out_387}=HA_cout_333+HA_out_334;
  assign {HA_cout_388,HA_out_388}=HA_cout_334+HA_out_335;
  assign {HA_cout_389,HA_out_389}=HA_cout_335+HA_out_336;
  assign {HA_cout_390,HA_out_390}=HA_cout_336+HA_out_337;
  assign {HA_cout_391,HA_out_391}=HA_cout_337+HA_out_338;
  assign {HA_cout_392,HA_out_392}=HA_cout_338+FA_out_3731;
  assign {HA_cout_393,HA_out_393}=FA_cout_3731+FA_out_3732;
  assign {HA_cout_394,HA_out_394}=FA_cout_3732+FA_out_3733;
  assign {HA_cout_395,HA_out_395}=FA_cout_3733+FA_out_3734;
  assign {HA_cout_396,HA_out_396}=FA_cout_3734+FA_out_3735;
  assign {HA_cout_397,HA_out_397}=FA_cout_3735+FA_out_3736;
  assign {HA_cout_398,HA_out_398}=FA_cout_3736+FA_out_3737;
  assign {HA_cout_399,HA_out_399}=FA_cout_3737+FA_out_3738;
  assign {HA_cout_400,HA_out_400}=FA_cout_3738+FA_out_3739;
  assign {HA_cout_401,HA_out_401}=FA_cout_3739+FA_out_3740;
  assign {HA_cout_402,HA_out_402}=FA_cout_3740+FA_out_3741;
  assign {HA_cout_403,HA_out_403}=FA_cout_3741+FA_out_3742;
  assign {HA_cout_404,HA_out_404}=FA_cout_3742+FA_out_3743;
  assign {HA_cout_405,HA_out_405}=FA_cout_3743+FA_out_3744;
  assign {HA_cout_406,HA_out_406}=FA_cout_3787+FA_out_3788;
  assign {HA_cout_407,HA_out_407}=FA_cout_3788+FA_out_3789;
  assign {HA_cout_408,HA_out_408}=FA_cout_3789+FA_out_3790;
  assign {HA_cout_409,HA_out_409}=FA_cout_3790+FA_out_3791;
  assign {HA_cout_410,HA_out_410}=FA_cout_3791+FA_out_3792;
  assign {HA_cout_411,HA_out_411}=FA_cout_3792+FA_out_3793;
  assign {HA_cout_412,HA_out_412}=FA_cout_3793+FA_out_3794;
  assign {HA_cout_413,HA_out_413}=FA_cout_3794+FA_out_3795;
  assign {HA_cout_414,HA_out_414}=FA_cout_3795+FA_out_3796;
  assign {HA_cout_415,HA_out_415}=FA_cout_3796+FA_out_3797;
  assign {HA_cout_416,HA_out_416}=FA_cout_3797+FA_out_3798;
  assign {HA_cout_417,HA_out_417}=FA_cout_3798+FA_out_3799;
  assign {HA_cout_418,HA_out_418}=FA_cout_3799+FA_out_3800;
  assign {HA_cout_419,HA_out_419}=FA_cout_3800+HA_out_341;
  assign {HA_cout_420,HA_out_420}=HA_cout_341+HA_out_342;
  assign {HA_cout_421,HA_out_421}=HA_cout_342+HA_out_343;
  assign {HA_cout_422,HA_out_422}=HA_cout_343+HA_out_344;
  assign {HA_cout_423,HA_out_423}=HA_cout_344+HA_out_345;
  assign {HA_cout_424,HA_out_424}=HA_cout_345+HA_out_346;
  assign {HA_cout_425,HA_out_425}=HA_cout_346+HA_out_347;
  assign {HA_cout_426,HA_out_426}=HA_cout_347+HA_out_348;
  assign {HA_cout_427,HA_out_427}=HA_cout_348+HA_out_349;
  assign {HA_cout_428,HA_out_428}=HA_cout_349+HA_out_350;
  assign {HA_cout_429,HA_out_429}=HA_cout_350+HA_out_351;
  assign {HA_cout_430,HA_out_430}=HA_cout_351+HA_out_352;
  assign {HA_cout_431,HA_out_431}=HA_cout_352+HA_out_353;
  assign {HA_cout_432,HA_out_432}=HA_cout_353+HA_out_354;
  assign {HA_cout_433,HA_out_433}=HA_cout_354+HA_out_355;
  assign {HA_cout_434,HA_out_434}=HA_cout_355+HA_out_356;
  assign {HA_cout_435,HA_out_435}=HA_cout_356+HA_out_357;
  assign {HA_cout_436,HA_out_436}=HA_cout_357+HA_out_358;
  assign {HA_cout_437,HA_out_437}=HA_cout_358+HA_out_359;
  assign {HA_cout_438,HA_out_438}=HA_cout_359+HA_out_360;
  assign {HA_cout_439,HA_out_439}=HA_cout_360+HA_out_361;
  assign {HA_cout_440,HA_out_440}=HA_cout_361+HA_out_362;
  assign {HA_cout_441,HA_out_441}=HA_cout_362+HA_out_363;
  assign {HA_cout_442,HA_out_442}=HA_cout_363+HA_out_364;
  assign {HA_cout_443,HA_out_443}=HA_cout_364+HA_out_365;
  assign {HA_cout_444,HA_out_444}=HA_cout_365+HA_out_366;
  assign {HA_cout_445,HA_out_445}=HA_cout_366+HA_out_367;
  assign {HA_cout_446,HA_out_446}=HA_cout_367+HA_out_368;
  assign {HA_cout_447,HA_out_447}=HA_cout_369+HA_out_370;
  assign {HA_cout_448,HA_out_448}=HA_cout_370+HA_out_371;
  assign {HA_cout_449,HA_out_449}=HA_cout_371+HA_out_372;
  assign {HA_cout_450,HA_out_450}=HA_cout_372+HA_out_373;
  assign {HA_cout_451,HA_out_451}=HA_cout_373+HA_out_374;
  assign {HA_cout_452,HA_out_452}=HA_cout_374+HA_out_375;
  assign {HA_cout_453,HA_out_453}=HA_cout_375+HA_out_376;
  assign {HA_cout_454,HA_out_454}=HA_cout_376+HA_out_377;
  assign {HA_cout_455,HA_out_455}=HA_cout_377+HA_out_378;
  assign {HA_cout_456,HA_out_456}=HA_cout_378+HA_out_379;
  assign {HA_cout_457,HA_out_457}=HA_cout_379+HA_out_380;
  assign {HA_cout_458,HA_out_458}=HA_cout_380+HA_out_381;
  assign {HA_cout_459,HA_out_459}=HA_cout_381+HA_out_382;
  assign {HA_cout_460,HA_out_460}=HA_cout_382+HA_out_383;
  assign {HA_cout_461,HA_out_461}=HA_cout_383+HA_out_384;
  assign {HA_cout_462,HA_out_462}=HA_cout_384+HA_out_385;
  assign {HA_cout_463,HA_out_463}=HA_cout_385+HA_out_386;
  assign {HA_cout_464,HA_out_464}=HA_cout_386+HA_out_387;
  assign {HA_cout_465,HA_out_465}=HA_cout_387+HA_out_388;
  assign {HA_cout_466,HA_out_466}=HA_cout_388+HA_out_389;
  assign {HA_cout_467,HA_out_467}=HA_cout_389+HA_out_390;
  assign {HA_cout_468,HA_out_468}=HA_cout_390+HA_out_391;
  assign {HA_cout_469,HA_out_469}=HA_cout_391+HA_out_392;
  assign {HA_cout_470,HA_out_470}=HA_cout_392+HA_out_393;
  assign {HA_cout_471,HA_out_471}=HA_cout_393+HA_out_394;
  assign {HA_cout_472,HA_out_472}=HA_cout_394+HA_out_395;
  assign {HA_cout_473,HA_out_473}=HA_cout_395+HA_out_396;
  assign {HA_cout_474,HA_out_474}=HA_cout_396+HA_out_397;
  assign {HA_cout_475,HA_out_475}=HA_cout_397+HA_out_398;
  assign {HA_cout_476,HA_out_476}=HA_cout_398+HA_out_399;
  assign {HA_cout_477,HA_out_477}=HA_cout_399+HA_out_400;
  assign {HA_cout_478,HA_out_478}=HA_cout_400+HA_out_401;
  assign {HA_cout_479,HA_out_479}=HA_cout_401+HA_out_402;
  assign {HA_cout_480,HA_out_480}=HA_cout_402+HA_out_403;
  assign {HA_cout_481,HA_out_481}=HA_cout_403+HA_out_404;
  assign {HA_cout_482,HA_out_482}=HA_cout_404+HA_out_405;
  assign {HA_cout_483,HA_out_483}=HA_cout_405+FA_out_3801;
  assign {HA_cout_484,HA_out_484}=FA_cout_3801+FA_out_3802;
  assign {HA_cout_485,HA_out_485}=FA_cout_3802+FA_out_3803;
  assign {HA_cout_486,HA_out_486}=FA_cout_3803+FA_out_3804;
  assign {HA_cout_487,HA_out_487}=FA_cout_3804+FA_out_3805;
  assign {HA_cout_488,HA_out_488}=FA_cout_3805+FA_out_3806;
  assign {HA_cout_489,HA_out_489}=FA_cout_3806+FA_out_3807;
  assign {HA_cout_490,HA_out_490}=FA_cout_3807+FA_out_3808;
  assign {HA_cout_491,HA_out_491}=FA_cout_3808+FA_out_3809;
  assign {HA_cout_492,HA_out_492}=FA_cout_3809+FA_out_3810;
  assign {HA_cout_493,HA_out_493}=FA_cout_3810+FA_out_3811;
  assign {HA_cout_494,HA_out_494}=FA_cout_3811+FA_out_3812;
  assign {HA_cout_495,HA_out_495}=FA_cout_3812+FA_out_3813;
  assign {HA_cout_496,HA_out_496}=FA_cout_3813+FA_out_3814;
  assign {HA_cout_497,HA_out_497}=FA_cout_3814+FA_out_3815;
  assign {HA_cout_498,HA_out_498}=FA_cout_3815+FA_out_3816;
  assign {HA_cout_499,HA_out_499}=FA_cout_3816+FA_out_3817;
  assign {HA_cout_500,HA_out_500}=FA_cout_3817+FA_out_3818;
  assign {HA_cout_501,HA_out_501}=FA_cout_3818+FA_out_3819;
  assign {HA_cout_502,HA_out_502}=FA_cout_3819+FA_out_3820;
  assign {HA_cout_503,HA_out_503}=FA_cout_3820+FA_out_3821;
  assign {HA_cout_504,HA_out_504}=FA_cout_3823+FA_out_3824;
  assign {HA_cout_505,HA_out_505}=FA_cout_3824+FA_out_3825;
  assign {HA_cout_506,HA_out_506}=FA_cout_3825+FA_out_3826;
  assign {HA_cout_507,HA_out_507}=FA_cout_3826+FA_out_3827;
  assign {HA_cout_508,HA_out_508}=FA_cout_3827+FA_out_3828;
  assign {HA_cout_509,HA_out_509}=FA_cout_3828+FA_out_3829;
  assign {HA_cout_510,HA_out_510}=FA_cout_3829+FA_out_3830;
  assign {HA_cout_511,HA_out_511}=FA_cout_3830+FA_out_3831;
  assign {HA_cout_512,HA_out_512}=FA_cout_3831+FA_out_3832;
  assign {HA_cout_513,HA_out_513}=FA_cout_3832+FA_out_3833;
  assign {HA_cout_514,HA_out_514}=FA_cout_3833+FA_out_3834;
  assign {HA_cout_515,HA_out_515}=FA_cout_3834+FA_out_3835;
  assign {HA_cout_516,HA_out_516}=FA_cout_3835+FA_out_3836;
  assign {HA_cout_517,HA_out_517}=FA_cout_3836+FA_out_3837;
  assign {HA_cout_518,HA_out_518}=FA_cout_3837+FA_out_3838;
  assign {HA_cout_519,HA_out_519}=FA_cout_3838+FA_out_3839;
  assign {HA_cout_520,HA_out_520}=FA_cout_3839+FA_out_3840;
  assign {HA_cout_521,HA_out_521}=FA_cout_3840+FA_out_3841;
  assign {HA_cout_522,HA_out_522}=FA_cout_3841+FA_out_3842;
  assign {HA_cout_523,HA_out_523}=FA_cout_3842+FA_out_3843;
  assign {HA_cout_524,HA_out_524}=FA_cout_3843+HA_out_406;
  assign {HA_cout_525,HA_out_525}=HA_cout_406+HA_out_407;
  assign {HA_cout_526,HA_out_526}=HA_cout_407+HA_out_408;
  assign {HA_cout_527,HA_out_527}=HA_cout_408+HA_out_409;
  assign {HA_cout_528,HA_out_528}=HA_cout_409+HA_out_410;
  assign {HA_cout_529,HA_out_529}=HA_cout_410+HA_out_411;
  assign {HA_cout_530,HA_out_530}=HA_cout_411+HA_out_412;
  assign {HA_cout_531,HA_out_531}=HA_cout_412+HA_out_413;
  assign {HA_cout_532,HA_out_532}=HA_cout_413+HA_out_414;
  assign {HA_cout_533,HA_out_533}=HA_cout_414+HA_out_415;
  assign {HA_cout_534,HA_out_534}=HA_cout_415+HA_out_416;
  assign {HA_cout_535,HA_out_535}=HA_cout_416+HA_out_417;
  assign {HA_cout_536,HA_out_536}=HA_cout_417+HA_out_418;
  assign {HA_cout_537,HA_out_537}=HA_cout_418+HA_out_419;
  assign {HA_cout_538,HA_out_538}=HA_cout_419+HA_out_420;
  assign {HA_cout_539,HA_out_539}=HA_cout_420+HA_out_421;
  assign {HA_cout_540,HA_out_540}=HA_cout_421+HA_out_422;
  assign {HA_cout_541,HA_out_541}=HA_cout_422+HA_out_423;
  assign {HA_cout_542,HA_out_542}=HA_cout_423+HA_out_424;
  assign {HA_cout_543,HA_out_543}=HA_cout_424+HA_out_425;
  assign {HA_cout_544,HA_out_544}=HA_cout_425+HA_out_426;
  assign {HA_cout_545,HA_out_545}=HA_cout_426+HA_out_427;
  assign {HA_cout_546,HA_out_546}=HA_cout_427+HA_out_428;
  assign {HA_cout_547,HA_out_547}=HA_cout_428+HA_out_429;
  assign {HA_cout_548,HA_out_548}=HA_cout_429+HA_out_430;
  assign {HA_cout_549,HA_out_549}=HA_cout_430+HA_out_431;
  assign {HA_cout_550,HA_out_550}=HA_cout_431+HA_out_432;
  assign {HA_cout_551,HA_out_551}=HA_cout_432+HA_out_433;
  assign {HA_cout_552,HA_out_552}=HA_cout_433+HA_out_434;
  assign {HA_cout_553,HA_out_553}=HA_cout_434+HA_out_435;
  assign {HA_cout_554,HA_out_554}=HA_cout_435+HA_out_436;
  assign {HA_cout_555,HA_out_555}=HA_cout_436+HA_out_437;
  assign {HA_cout_556,HA_out_556}=HA_cout_437+HA_out_438;
  assign {HA_cout_557,HA_out_557}=HA_cout_438+HA_out_439;
  assign {HA_cout_558,HA_out_558}=HA_cout_439+HA_out_440;
  assign {HA_cout_559,HA_out_559}=HA_cout_440+HA_out_441;
  assign {HA_cout_560,HA_out_560}=HA_cout_441+HA_out_442;
  assign {HA_cout_561,HA_out_561}=HA_cout_442+HA_out_443;
  assign {HA_cout_562,HA_out_562}=HA_cout_443+HA_out_444;
  assign {HA_cout_563,HA_out_563}=HA_cout_444+HA_out_445;
  assign {HA_cout_564,HA_out_564}=HA_cout_445+HA_out_446;
  assign {HA_cout_565,HA_out_565}=HA_cout_446+HA_cout_368;


  always @(*)
  begin
      REGS_0<=inp_0[0];
      REGS_1<=HA_out_0;
      REGS_2<=HA_out_42;
      REGS_3<=HA_cout_42;
      REGS_4<=FA_cout_1323;
      REGS_5<=FA_cout_1324;
      REGS_6<=FA_cout_1325;
      REGS_7<=FA_cout_1326;
      REGS_8<=FA_cout_1327;
      REGS_9<=FA_cout_1328;
      REGS_10<=FA_cout_1329;
      REGS_11<=FA_cout_1330;
      REGS_12<=FA_cout_1331;
      REGS_13<=FA_cout_1332;
      REGS_14<=FA_cout_1333;
      REGS_15<=FA_cout_1334;
      REGS_16<=FA_cout_1335;
      REGS_17<=FA_cout_1336;
      REGS_18<=FA_cout_1337;
      REGS_19<=FA_cout_1338;
      REGS_20<=FA_cout_1339;
      REGS_21<=FA_cout_1340;
      REGS_22<=FA_cout_1341;
      REGS_23<=FA_cout_1342;
      REGS_24<=FA_cout_1343;
      REGS_25<=FA_cout_1344;
      REGS_26<=FA_cout_1345;
      REGS_27<=FA_cout_1346;
      REGS_28<=FA_cout_1347;
      REGS_29<=FA_cout_1348;
      REGS_30<=FA_cout_1349;
      REGS_31<=FA_cout_1350;
      REGS_32<=FA_cout_1351;
      REGS_33<=FA_cout_1352;
      REGS_34<=FA_cout_1353;
      REGS_35<=FA_cout_1354;
      REGS_36<=FA_cout_1355;
      REGS_37<=FA_cout_1356;
      REGS_38<=FA_cout_1357;
      REGS_39<=FA_cout_1358;
      REGS_40<=FA_cout_1359;
      REGS_41<=FA_cout_1360;
      REGS_42<=FA_cout_1361;
      REGS_43<=FA_cout_1362;
      REGS_44<=FA_cout_1363;
      REGS_45<=FA_cout_1364;
      REGS_46<=FA_cout_1365;
      REGS_47<=FA_cout_1366;
      REGS_48<=FA_cout_1367;
      REGS_49<=FA_cout_1368;
      REGS_50<=FA_cout_1369;
      REGS_51<=FA_cout_1370;
      REGS_52<=FA_cout_1371;
      REGS_53<=FA_cout_1372;
      REGS_54<=FA_cout_1373;
      REGS_55<=FA_cout_1374;
      REGS_56<=FA_cout_1375;
      REGS_57<=FA_cout_1376;
      REGS_58<=FA_cout_1377;
      REGS_59<=FA_cout_1378;
      REGS_60<=FA_cout_1379;
      REGS_61<=FA_cout_1380;
      REGS_62<=FA_cout_1381;
      REGS_63<=FA_cout_1382;
      REGS_64<=FA_cout_1383;
      REGS_65<=FA_cout_1384;
      REGS_66<=FA_cout_1385;
      REGS_67<=FA_out_1323;
      REGS_68<=FA_out_1324;
      REGS_69<=FA_out_1325;
      REGS_70<=FA_out_1326;
      REGS_71<=FA_out_1327;
      REGS_72<=FA_out_1328;
      REGS_73<=FA_out_1329;
      REGS_74<=FA_out_1330;
      REGS_75<=FA_out_1331;
      REGS_76<=FA_out_1332;
      REGS_77<=FA_out_1333;
      REGS_78<=FA_out_1334;
      REGS_79<=FA_out_1335;
      REGS_80<=FA_out_1336;
      REGS_81<=FA_out_1337;
      REGS_82<=FA_out_1338;
      REGS_83<=FA_out_1339;
      REGS_84<=FA_out_1340;
      REGS_85<=FA_out_1341;
      REGS_86<=FA_out_1342;
      REGS_87<=FA_out_1343;
      REGS_88<=FA_out_1344;
      REGS_89<=FA_out_1345;
      REGS_90<=FA_out_1346;
      REGS_91<=FA_out_1347;
      REGS_92<=FA_out_1348;
      REGS_93<=FA_out_1349;
      REGS_94<=FA_out_1350;
      REGS_95<=FA_out_1351;
      REGS_96<=FA_out_1352;
      REGS_97<=FA_out_1353;
      REGS_98<=FA_out_1354;
      REGS_99<=FA_out_1355;
      REGS_100<=FA_out_1356;
      REGS_101<=FA_out_1357;
      REGS_102<=FA_out_1358;
      REGS_103<=FA_out_1359;
      REGS_104<=FA_out_1360;
      REGS_105<=FA_out_1361;
      REGS_106<=FA_out_1362;
      REGS_107<=FA_out_1363;
      REGS_108<=FA_out_1364;
      REGS_109<=FA_out_1365;
      REGS_110<=FA_out_1366;
      REGS_111<=FA_out_1367;
      REGS_112<=FA_out_1368;
      REGS_113<=FA_out_1369;
      REGS_114<=FA_out_1370;
      REGS_115<=FA_out_1371;
      REGS_116<=FA_out_1372;
      REGS_117<=FA_out_1373;
      REGS_118<=FA_out_1374;
      REGS_119<=FA_out_1375;
      REGS_120<=FA_out_1376;
      REGS_121<=FA_out_1377;
      REGS_122<=FA_out_1378;
      REGS_123<=FA_out_1379;
      REGS_124<=FA_out_1380;
      REGS_125<=FA_out_1381;
      REGS_126<=FA_out_1382;
      REGS_127<=FA_out_1383;
      REGS_128<=FA_out_1384;
      REGS_129<=FA_out_1385;
      REGS_130<=FA_out_1386;
      REGS_131<=FA_cout_1386;
      REGS_132<=FA_out_1387;
      REGS_133<=FA_cout_1387;
      REGS_134<=FA_out_64;
      REGS_135<=HA_out_43;
      REGS_136<=HA_cout_43;
      REGS_137<=HA_cout_44;
      REGS_138<=FA_cout_1388;
      REGS_139<=FA_cout_1389;
      REGS_140<=FA_cout_1390;
      REGS_141<=FA_cout_1391;
      REGS_142<=FA_cout_1392;
      REGS_143<=FA_cout_1393;
      REGS_144<=FA_cout_1394;
      REGS_145<=FA_cout_1395;
      REGS_146<=FA_cout_1396;
      REGS_147<=FA_cout_1397;
      REGS_148<=FA_cout_1398;
      REGS_149<=FA_cout_1399;
      REGS_150<=FA_cout_1400;
      REGS_151<=FA_cout_1401;
      REGS_152<=FA_cout_1402;
      REGS_153<=FA_cout_1403;
      REGS_154<=FA_cout_1404;
      REGS_155<=FA_cout_1405;
      REGS_156<=FA_cout_1406;
      REGS_157<=FA_cout_1407;
      REGS_158<=FA_cout_1408;
      REGS_159<=FA_cout_1409;
      REGS_160<=FA_cout_1410;
      REGS_161<=FA_cout_1411;
      REGS_162<=FA_cout_1412;
      REGS_163<=FA_cout_1413;
      REGS_164<=FA_cout_1414;
      REGS_165<=FA_cout_1415;
      REGS_166<=FA_cout_1416;
      REGS_167<=FA_cout_1417;
      REGS_168<=FA_cout_1418;
      REGS_169<=FA_cout_1419;
      REGS_170<=FA_cout_1420;
      REGS_171<=FA_cout_1421;
      REGS_172<=FA_cout_1422;
      REGS_173<=FA_cout_1423;
      REGS_174<=FA_cout_1424;
      REGS_175<=FA_cout_1425;
      REGS_176<=FA_cout_1426;
      REGS_177<=FA_cout_1427;
      REGS_178<=FA_cout_1428;
      REGS_179<=FA_cout_1429;
      REGS_180<=FA_cout_1430;
      REGS_181<=FA_cout_1431;
      REGS_182<=FA_cout_1432;
      REGS_183<=FA_cout_1433;
      REGS_184<=FA_cout_1434;
      REGS_185<=FA_cout_1435;
      REGS_186<=FA_cout_1436;
      REGS_187<=FA_cout_1437;
      REGS_188<=FA_cout_1438;
      REGS_189<=FA_cout_1439;
      REGS_190<=FA_cout_1440;
      REGS_191<=FA_cout_1441;
      REGS_192<=FA_cout_1442;
      REGS_193<=FA_cout_1443;
      REGS_194<=FA_cout_1444;
      REGS_195<=FA_out_1445;
      REGS_196<=FA_cout_1445;
      REGS_197<=HA_out_44;
      REGS_198<=FA_out_1388;
      REGS_199<=FA_out_1389;
      REGS_200<=FA_out_1390;
      REGS_201<=FA_out_1391;
      REGS_202<=FA_out_1392;
      REGS_203<=FA_out_1393;
      REGS_204<=FA_out_1394;
      REGS_205<=FA_out_1395;
      REGS_206<=FA_out_1396;
      REGS_207<=FA_out_1397;
      REGS_208<=FA_out_1398;
      REGS_209<=FA_out_1399;
      REGS_210<=FA_out_1400;
      REGS_211<=FA_out_1401;
      REGS_212<=FA_out_1402;
      REGS_213<=FA_out_1403;
      REGS_214<=FA_out_1404;
      REGS_215<=FA_out_1405;
      REGS_216<=FA_out_1406;
      REGS_217<=FA_out_1407;
      REGS_218<=FA_out_1408;
      REGS_219<=FA_out_1409;
      REGS_220<=FA_out_1410;
      REGS_221<=FA_out_1411;
      REGS_222<=FA_out_1412;
      REGS_223<=FA_out_1413;
      REGS_224<=FA_out_1414;
      REGS_225<=FA_out_1415;
      REGS_226<=FA_out_1416;
      REGS_227<=FA_out_1417;
      REGS_228<=FA_out_1418;
      REGS_229<=FA_out_1419;
      REGS_230<=FA_out_1420;
      REGS_231<=FA_out_1421;
      REGS_232<=FA_out_1422;
      REGS_233<=FA_out_1423;
      REGS_234<=FA_out_1424;
      REGS_235<=FA_out_1425;
      REGS_236<=FA_out_1426;
      REGS_237<=FA_out_1427;
      REGS_238<=FA_out_1428;
      REGS_239<=FA_out_1429;
      REGS_240<=FA_out_1430;
      REGS_241<=FA_out_1431;
      REGS_242<=FA_out_1432;
      REGS_243<=FA_out_1433;
      REGS_244<=FA_out_1434;
      REGS_245<=FA_out_1435;
      REGS_246<=FA_out_1436;
      REGS_247<=FA_out_1437;
      REGS_248<=FA_out_1438;
      REGS_249<=FA_out_1439;
      REGS_250<=FA_out_1440;
      REGS_251<=FA_out_1441;
      REGS_252<=FA_out_1442;
      REGS_253<=FA_out_1443;
      REGS_254<=FA_out_1444;
      REGS_255<=FA_out_1446;
      REGS_256<=FA_cout_1446;
      REGS_257<=FA_out_1447;
      REGS_258<=FA_cout_1447;
      REGS_259<=FA_out_1448;
      REGS_260<=FA_cout_1448;
      REGS_261<=FA_out_1449;
      REGS_262<=FA_cout_1449;
      REGS_263<=FA_out_1450;
      REGS_264<=FA_cout_1450;
      REGS_265<=FA_out_1451;
      REGS_266<=FA_cout_1451;
      REGS_267<=FA_out_1452;
      REGS_268<=FA_cout_1452;
      REGS_269<=FA_out_1453;
      REGS_270<=FA_cout_1453;
      REGS_271<=inp_9[0];
      REGS_272<=HA_out_3;
      REGS_273<=HA_out_45;
      REGS_274<=HA_cout_45;
      REGS_275<=FA_cout_1454;
      REGS_276<=FA_cout_1455;
      REGS_277<=FA_cout_1456;
      REGS_278<=FA_cout_1457;
      REGS_279<=FA_cout_1458;
      REGS_280<=FA_cout_1459;
      REGS_281<=FA_cout_1460;
      REGS_282<=FA_cout_1461;
      REGS_283<=FA_cout_1462;
      REGS_284<=FA_cout_1463;
      REGS_285<=FA_cout_1464;
      REGS_286<=FA_cout_1465;
      REGS_287<=FA_cout_1466;
      REGS_288<=FA_cout_1467;
      REGS_289<=FA_cout_1468;
      REGS_290<=FA_cout_1469;
      REGS_291<=FA_cout_1470;
      REGS_292<=FA_cout_1471;
      REGS_293<=FA_cout_1472;
      REGS_294<=FA_cout_1473;
      REGS_295<=FA_cout_1474;
      REGS_296<=FA_cout_1475;
      REGS_297<=FA_cout_1476;
      REGS_298<=FA_cout_1477;
      REGS_299<=FA_cout_1478;
      REGS_300<=FA_cout_1479;
      REGS_301<=FA_cout_1480;
      REGS_302<=FA_cout_1481;
      REGS_303<=FA_cout_1482;
      REGS_304<=FA_cout_1483;
      REGS_305<=FA_cout_1484;
      REGS_306<=FA_cout_1485;
      REGS_307<=FA_cout_1486;
      REGS_308<=FA_cout_1487;
      REGS_309<=FA_cout_1488;
      REGS_310<=FA_cout_1489;
      REGS_311<=FA_cout_1490;
      REGS_312<=FA_cout_1491;
      REGS_313<=FA_cout_1492;
      REGS_314<=FA_cout_1493;
      REGS_315<=FA_cout_1494;
      REGS_316<=FA_cout_1495;
      REGS_317<=FA_cout_1496;
      REGS_318<=FA_cout_1497;
      REGS_319<=FA_cout_1498;
      REGS_320<=FA_cout_1499;
      REGS_321<=FA_cout_1500;
      REGS_322<=FA_cout_1501;
      REGS_323<=FA_cout_1502;
      REGS_324<=FA_cout_1503;
      REGS_325<=FA_cout_1504;
      REGS_326<=FA_cout_1505;
      REGS_327<=FA_cout_1506;
      REGS_328<=FA_cout_1507;
      REGS_329<=FA_out_1508;
      REGS_330<=FA_cout_1508;
      REGS_331<=FA_out_1509;
      REGS_332<=FA_cout_1509;
      REGS_333<=FA_out_1454;
      REGS_334<=FA_out_1455;
      REGS_335<=FA_out_1456;
      REGS_336<=FA_out_1457;
      REGS_337<=FA_out_1458;
      REGS_338<=FA_out_1459;
      REGS_339<=FA_out_1460;
      REGS_340<=FA_out_1461;
      REGS_341<=FA_out_1462;
      REGS_342<=FA_out_1463;
      REGS_343<=FA_out_1464;
      REGS_344<=FA_out_1465;
      REGS_345<=FA_out_1466;
      REGS_346<=FA_out_1467;
      REGS_347<=FA_out_1468;
      REGS_348<=FA_out_1469;
      REGS_349<=FA_out_1470;
      REGS_350<=FA_out_1471;
      REGS_351<=FA_out_1472;
      REGS_352<=FA_out_1473;
      REGS_353<=FA_out_1474;
      REGS_354<=FA_out_1475;
      REGS_355<=FA_out_1476;
      REGS_356<=FA_out_1477;
      REGS_357<=FA_out_1478;
      REGS_358<=FA_out_1479;
      REGS_359<=FA_out_1480;
      REGS_360<=FA_out_1481;
      REGS_361<=FA_out_1482;
      REGS_362<=FA_out_1483;
      REGS_363<=FA_out_1484;
      REGS_364<=FA_out_1485;
      REGS_365<=FA_out_1486;
      REGS_366<=FA_out_1487;
      REGS_367<=FA_out_1488;
      REGS_368<=FA_out_1489;
      REGS_369<=FA_out_1490;
      REGS_370<=FA_out_1491;
      REGS_371<=FA_out_1492;
      REGS_372<=FA_out_1493;
      REGS_373<=FA_out_1494;
      REGS_374<=FA_out_1495;
      REGS_375<=FA_out_1496;
      REGS_376<=FA_out_1497;
      REGS_377<=FA_out_1498;
      REGS_378<=FA_out_1499;
      REGS_379<=FA_out_1500;
      REGS_380<=FA_out_1501;
      REGS_381<=FA_out_1502;
      REGS_382<=FA_out_1503;
      REGS_383<=FA_out_1504;
      REGS_384<=FA_out_1505;
      REGS_385<=FA_out_1506;
      REGS_386<=FA_out_1507;
      REGS_387<=FA_out_1510;
      REGS_388<=FA_cout_1510;
      REGS_389<=FA_out_1511;
      REGS_390<=FA_cout_1511;
      REGS_391<=FA_out_1512;
      REGS_392<=FA_cout_1512;
      REGS_393<=FA_out_1513;
      REGS_394<=FA_cout_1513;
      REGS_395<=FA_out_1514;
      REGS_396<=FA_cout_1514;
      REGS_397<=FA_out_1515;
      REGS_398<=FA_cout_1515;
      REGS_399<=FA_out_1516;
      REGS_400<=FA_cout_1516;
      REGS_401<=FA_out_1517;
      REGS_402<=FA_cout_1517;
      REGS_403<=FA_out_256;
      REGS_404<=HA_out_46;
      REGS_405<=HA_cout_46;
      REGS_406<=HA_cout_47;
      REGS_407<=FA_cout_1518;
      REGS_408<=FA_cout_1519;
      REGS_409<=FA_cout_1520;
      REGS_410<=FA_cout_1521;
      REGS_411<=FA_cout_1522;
      REGS_412<=FA_cout_1523;
      REGS_413<=FA_cout_1524;
      REGS_414<=FA_cout_1525;
      REGS_415<=FA_cout_1526;
      REGS_416<=FA_cout_1527;
      REGS_417<=FA_cout_1528;
      REGS_418<=FA_cout_1529;
      REGS_419<=FA_cout_1530;
      REGS_420<=FA_cout_1531;
      REGS_421<=FA_cout_1532;
      REGS_422<=FA_cout_1533;
      REGS_423<=FA_cout_1534;
      REGS_424<=FA_cout_1535;
      REGS_425<=FA_cout_1536;
      REGS_426<=FA_cout_1537;
      REGS_427<=FA_cout_1538;
      REGS_428<=FA_cout_1539;
      REGS_429<=FA_cout_1540;
      REGS_430<=FA_cout_1541;
      REGS_431<=FA_cout_1542;
      REGS_432<=FA_cout_1543;
      REGS_433<=FA_cout_1544;
      REGS_434<=FA_cout_1545;
      REGS_435<=FA_cout_1546;
      REGS_436<=FA_cout_1547;
      REGS_437<=FA_cout_1548;
      REGS_438<=FA_cout_1549;
      REGS_439<=FA_cout_1550;
      REGS_440<=FA_cout_1551;
      REGS_441<=FA_cout_1552;
      REGS_442<=FA_cout_1553;
      REGS_443<=FA_cout_1554;
      REGS_444<=FA_cout_1555;
      REGS_445<=FA_cout_1556;
      REGS_446<=FA_cout_1557;
      REGS_447<=FA_cout_1558;
      REGS_448<=FA_cout_1559;
      REGS_449<=FA_cout_1560;
      REGS_450<=FA_cout_1561;
      REGS_451<=FA_cout_1562;
      REGS_452<=FA_cout_1563;
      REGS_453<=FA_cout_1564;
      REGS_454<=FA_cout_1565;
      REGS_455<=FA_out_1566;
      REGS_456<=FA_cout_1566;
      REGS_457<=FA_out_1567;
      REGS_458<=FA_cout_1567;
      REGS_459<=FA_out_1568;
      REGS_460<=FA_cout_1568;
      REGS_461<=HA_out_47;
      REGS_462<=FA_out_1518;
      REGS_463<=FA_out_1519;
      REGS_464<=FA_out_1520;
      REGS_465<=FA_out_1521;
      REGS_466<=FA_out_1522;
      REGS_467<=FA_out_1523;
      REGS_468<=FA_out_1524;
      REGS_469<=FA_out_1525;
      REGS_470<=FA_out_1526;
      REGS_471<=FA_out_1527;
      REGS_472<=FA_out_1528;
      REGS_473<=FA_out_1529;
      REGS_474<=FA_out_1530;
      REGS_475<=FA_out_1531;
      REGS_476<=FA_out_1532;
      REGS_477<=FA_out_1533;
      REGS_478<=FA_out_1534;
      REGS_479<=FA_out_1535;
      REGS_480<=FA_out_1536;
      REGS_481<=FA_out_1537;
      REGS_482<=FA_out_1538;
      REGS_483<=FA_out_1539;
      REGS_484<=FA_out_1540;
      REGS_485<=FA_out_1541;
      REGS_486<=FA_out_1542;
      REGS_487<=FA_out_1543;
      REGS_488<=FA_out_1544;
      REGS_489<=FA_out_1545;
      REGS_490<=FA_out_1546;
      REGS_491<=FA_out_1547;
      REGS_492<=FA_out_1548;
      REGS_493<=FA_out_1549;
      REGS_494<=FA_out_1550;
      REGS_495<=FA_out_1551;
      REGS_496<=FA_out_1552;
      REGS_497<=FA_out_1553;
      REGS_498<=FA_out_1554;
      REGS_499<=FA_out_1555;
      REGS_500<=FA_out_1556;
      REGS_501<=FA_out_1557;
      REGS_502<=FA_out_1558;
      REGS_503<=FA_out_1559;
      REGS_504<=FA_out_1560;
      REGS_505<=FA_out_1561;
      REGS_506<=FA_out_1562;
      REGS_507<=FA_out_1563;
      REGS_508<=FA_out_1564;
      REGS_509<=FA_out_1565;
      REGS_510<=FA_out_1569;
      REGS_511<=FA_cout_1569;
      REGS_512<=FA_out_1570;
      REGS_513<=FA_cout_1570;
      REGS_514<=FA_out_1571;
      REGS_515<=FA_cout_1571;
      REGS_516<=FA_out_1572;
      REGS_517<=FA_cout_1572;
      REGS_518<=FA_out_1573;
      REGS_519<=FA_cout_1573;
      REGS_520<=FA_out_1574;
      REGS_521<=FA_cout_1574;
      REGS_522<=FA_out_1575;
      REGS_523<=FA_cout_1575;
      REGS_524<=FA_out_1576;
      REGS_525<=FA_cout_1576;
      REGS_526<=FA_out_1577;
      REGS_527<=FA_cout_1577;
      REGS_528<=FA_out_1578;
      REGS_529<=FA_cout_1578;
      REGS_530<=FA_out_1579;
      REGS_531<=FA_cout_1579;
      REGS_532<=FA_out_1580;
      REGS_533<=FA_cout_1580;
      REGS_534<=FA_out_1581;
      REGS_535<=FA_cout_1581;
      REGS_536<=FA_out_1582;
      REGS_537<=FA_cout_1582;
      REGS_538<=FA_out_1583;
      REGS_539<=FA_cout_1583;
      REGS_540<=FA_out_1584;
      REGS_541<=FA_cout_1584;
      REGS_542<=inp_18[0];
      REGS_543<=HA_out_6;
      REGS_544<=HA_out_48;
      REGS_545<=HA_cout_48;
      REGS_546<=FA_cout_1585;
      REGS_547<=FA_cout_1586;
      REGS_548<=FA_cout_1587;
      REGS_549<=FA_cout_1588;
      REGS_550<=FA_cout_1589;
      REGS_551<=FA_cout_1590;
      REGS_552<=FA_cout_1591;
      REGS_553<=FA_cout_1592;
      REGS_554<=FA_cout_1593;
      REGS_555<=FA_cout_1594;
      REGS_556<=FA_cout_1595;
      REGS_557<=FA_cout_1596;
      REGS_558<=FA_cout_1597;
      REGS_559<=FA_cout_1598;
      REGS_560<=FA_cout_1599;
      REGS_561<=FA_cout_1600;
      REGS_562<=FA_cout_1601;
      REGS_563<=FA_cout_1602;
      REGS_564<=FA_cout_1603;
      REGS_565<=FA_cout_1604;
      REGS_566<=FA_cout_1605;
      REGS_567<=FA_cout_1606;
      REGS_568<=FA_cout_1607;
      REGS_569<=FA_cout_1608;
      REGS_570<=FA_cout_1609;
      REGS_571<=FA_cout_1610;
      REGS_572<=FA_cout_1611;
      REGS_573<=FA_cout_1612;
      REGS_574<=FA_cout_1613;
      REGS_575<=FA_cout_1614;
      REGS_576<=FA_cout_1615;
      REGS_577<=FA_cout_1616;
      REGS_578<=FA_cout_1617;
      REGS_579<=FA_cout_1618;
      REGS_580<=FA_cout_1619;
      REGS_581<=FA_cout_1620;
      REGS_582<=FA_cout_1621;
      REGS_583<=FA_cout_1622;
      REGS_584<=FA_cout_1623;
      REGS_585<=FA_cout_1624;
      REGS_586<=FA_cout_1625;
      REGS_587<=FA_cout_1626;
      REGS_588<=FA_cout_1627;
      REGS_589<=FA_cout_1628;
      REGS_590<=FA_cout_1629;
      REGS_591<=FA_out_1630;
      REGS_592<=FA_cout_1630;
      REGS_593<=FA_out_1631;
      REGS_594<=FA_cout_1631;
      REGS_595<=FA_out_1632;
      REGS_596<=FA_cout_1632;
      REGS_597<=FA_out_1633;
      REGS_598<=FA_cout_1633;
      REGS_599<=FA_out_1585;
      REGS_600<=FA_out_1586;
      REGS_601<=FA_out_1587;
      REGS_602<=FA_out_1588;
      REGS_603<=FA_out_1589;
      REGS_604<=FA_out_1590;
      REGS_605<=FA_out_1591;
      REGS_606<=FA_out_1592;
      REGS_607<=FA_out_1593;
      REGS_608<=FA_out_1594;
      REGS_609<=FA_out_1595;
      REGS_610<=FA_out_1596;
      REGS_611<=FA_out_1597;
      REGS_612<=FA_out_1598;
      REGS_613<=FA_out_1599;
      REGS_614<=FA_out_1600;
      REGS_615<=FA_out_1601;
      REGS_616<=FA_out_1602;
      REGS_617<=FA_out_1603;
      REGS_618<=FA_out_1604;
      REGS_619<=FA_out_1605;
      REGS_620<=FA_out_1606;
      REGS_621<=FA_out_1607;
      REGS_622<=FA_out_1608;
      REGS_623<=FA_out_1609;
      REGS_624<=FA_out_1610;
      REGS_625<=FA_out_1611;
      REGS_626<=FA_out_1612;
      REGS_627<=FA_out_1613;
      REGS_628<=FA_out_1614;
      REGS_629<=FA_out_1615;
      REGS_630<=FA_out_1616;
      REGS_631<=FA_out_1617;
      REGS_632<=FA_out_1618;
      REGS_633<=FA_out_1619;
      REGS_634<=FA_out_1620;
      REGS_635<=FA_out_1621;
      REGS_636<=FA_out_1622;
      REGS_637<=FA_out_1623;
      REGS_638<=FA_out_1624;
      REGS_639<=FA_out_1625;
      REGS_640<=FA_out_1626;
      REGS_641<=FA_out_1627;
      REGS_642<=FA_out_1628;
      REGS_643<=FA_out_1629;
      REGS_644<=FA_out_1634;
      REGS_645<=FA_cout_1634;
      REGS_646<=FA_out_1635;
      REGS_647<=FA_cout_1635;
      REGS_648<=FA_out_1636;
      REGS_649<=FA_cout_1636;
      REGS_650<=FA_out_1637;
      REGS_651<=FA_cout_1637;
      REGS_652<=FA_out_1638;
      REGS_653<=FA_cout_1638;
      REGS_654<=FA_out_1639;
      REGS_655<=FA_cout_1639;
      REGS_656<=FA_out_1640;
      REGS_657<=FA_cout_1640;
      REGS_658<=FA_out_1641;
      REGS_659<=FA_cout_1641;
      REGS_660<=FA_out_1642;
      REGS_661<=FA_cout_1642;
      REGS_662<=FA_out_1643;
      REGS_663<=FA_cout_1643;
      REGS_664<=FA_out_1644;
      REGS_665<=FA_cout_1644;
      REGS_666<=FA_out_1645;
      REGS_667<=FA_cout_1645;
      REGS_668<=FA_out_1646;
      REGS_669<=FA_cout_1646;
      REGS_670<=FA_out_1647;
      REGS_671<=FA_cout_1647;
      REGS_672<=FA_out_448;
      REGS_673<=HA_out_49;
      REGS_674<=HA_cout_49;
      REGS_675<=HA_cout_50;
      REGS_676<=FA_cout_1648;
      REGS_677<=FA_cout_1649;
      REGS_678<=FA_cout_1650;
      REGS_679<=FA_cout_1651;
      REGS_680<=FA_cout_1652;
      REGS_681<=FA_cout_1653;
      REGS_682<=FA_cout_1654;
      REGS_683<=FA_cout_1655;
      REGS_684<=FA_cout_1656;
      REGS_685<=FA_cout_1657;
      REGS_686<=FA_cout_1658;
      REGS_687<=FA_cout_1659;
      REGS_688<=FA_cout_1660;
      REGS_689<=FA_cout_1661;
      REGS_690<=FA_cout_1662;
      REGS_691<=FA_cout_1663;
      REGS_692<=FA_cout_1664;
      REGS_693<=FA_cout_1665;
      REGS_694<=FA_cout_1666;
      REGS_695<=FA_cout_1667;
      REGS_696<=FA_cout_1668;
      REGS_697<=FA_cout_1669;
      REGS_698<=FA_cout_1670;
      REGS_699<=FA_cout_1671;
      REGS_700<=FA_cout_1672;
      REGS_701<=FA_cout_1673;
      REGS_702<=FA_cout_1674;
      REGS_703<=FA_cout_1675;
      REGS_704<=FA_cout_1676;
      REGS_705<=FA_cout_1677;
      REGS_706<=FA_cout_1678;
      REGS_707<=FA_cout_1679;
      REGS_708<=FA_cout_1680;
      REGS_709<=FA_cout_1681;
      REGS_710<=FA_cout_1682;
      REGS_711<=FA_cout_1683;
      REGS_712<=FA_cout_1684;
      REGS_713<=FA_cout_1685;
      REGS_714<=FA_cout_1686;
      REGS_715<=FA_out_1687;
      REGS_716<=FA_cout_1687;
      REGS_717<=FA_out_1688;
      REGS_718<=FA_cout_1688;
      REGS_719<=FA_out_1689;
      REGS_720<=FA_cout_1689;
      REGS_721<=FA_out_1690;
      REGS_722<=FA_cout_1690;
      REGS_723<=FA_out_1691;
      REGS_724<=FA_cout_1691;
      REGS_725<=HA_out_50;
      REGS_726<=FA_out_1648;
      REGS_727<=FA_out_1649;
      REGS_728<=FA_out_1650;
      REGS_729<=FA_out_1651;
      REGS_730<=FA_out_1652;
      REGS_731<=FA_out_1653;
      REGS_732<=FA_out_1654;
      REGS_733<=FA_out_1655;
      REGS_734<=FA_out_1656;
      REGS_735<=FA_out_1657;
      REGS_736<=FA_out_1658;
      REGS_737<=FA_out_1659;
      REGS_738<=FA_out_1660;
      REGS_739<=FA_out_1661;
      REGS_740<=FA_out_1662;
      REGS_741<=FA_out_1663;
      REGS_742<=FA_out_1664;
      REGS_743<=FA_out_1665;
      REGS_744<=FA_out_1666;
      REGS_745<=FA_out_1667;
      REGS_746<=FA_out_1668;
      REGS_747<=FA_out_1669;
      REGS_748<=FA_out_1670;
      REGS_749<=FA_out_1671;
      REGS_750<=FA_out_1672;
      REGS_751<=FA_out_1673;
      REGS_752<=FA_out_1674;
      REGS_753<=FA_out_1675;
      REGS_754<=FA_out_1676;
      REGS_755<=FA_out_1677;
      REGS_756<=FA_out_1678;
      REGS_757<=FA_out_1679;
      REGS_758<=FA_out_1680;
      REGS_759<=FA_out_1681;
      REGS_760<=FA_out_1682;
      REGS_761<=FA_out_1683;
      REGS_762<=FA_out_1684;
      REGS_763<=FA_out_1685;
      REGS_764<=FA_out_1686;
      REGS_765<=FA_out_1692;
      REGS_766<=FA_cout_1692;
      REGS_767<=FA_out_1693;
      REGS_768<=FA_cout_1693;
      REGS_769<=FA_out_1694;
      REGS_770<=FA_cout_1694;
      REGS_771<=FA_out_1695;
      REGS_772<=FA_cout_1695;
      REGS_773<=FA_out_1696;
      REGS_774<=FA_cout_1696;
      REGS_775<=FA_out_1697;
      REGS_776<=FA_cout_1697;
      REGS_777<=FA_out_1698;
      REGS_778<=FA_cout_1698;
      REGS_779<=FA_out_1699;
      REGS_780<=FA_cout_1699;
      REGS_781<=FA_out_1700;
      REGS_782<=FA_cout_1700;
      REGS_783<=FA_out_1701;
      REGS_784<=FA_cout_1701;
      REGS_785<=FA_out_1702;
      REGS_786<=FA_cout_1702;
      REGS_787<=FA_out_1703;
      REGS_788<=FA_cout_1703;
      REGS_789<=FA_out_1704;
      REGS_790<=FA_cout_1704;
      REGS_791<=FA_out_1705;
      REGS_792<=FA_cout_1705;
      REGS_793<=FA_out_1706;
      REGS_794<=FA_cout_1706;
      REGS_795<=FA_out_1707;
      REGS_796<=FA_cout_1707;
      REGS_797<=FA_out_1708;
      REGS_798<=FA_cout_1708;
      REGS_799<=FA_out_1709;
      REGS_800<=FA_cout_1709;
      REGS_801<=FA_out_1710;
      REGS_802<=FA_cout_1710;
      REGS_803<=FA_out_1711;
      REGS_804<=FA_cout_1711;
      REGS_805<=FA_out_1712;
      REGS_806<=FA_cout_1712;
      REGS_807<=FA_out_1713;
      REGS_808<=FA_cout_1713;
      REGS_809<=FA_out_1714;
      REGS_810<=FA_cout_1714;
      REGS_811<=FA_out_1715;
      REGS_812<=FA_cout_1715;
      REGS_813<=inp_27[0];
      REGS_814<=HA_out_9;
      REGS_815<=HA_out_51;
      REGS_816<=HA_cout_51;
      REGS_817<=FA_cout_1716;
      REGS_818<=FA_cout_1717;
      REGS_819<=FA_cout_1718;
      REGS_820<=FA_cout_1719;
      REGS_821<=FA_cout_1720;
      REGS_822<=FA_cout_1721;
      REGS_823<=FA_cout_1722;
      REGS_824<=FA_cout_1723;
      REGS_825<=FA_cout_1724;
      REGS_826<=FA_cout_1725;
      REGS_827<=FA_cout_1726;
      REGS_828<=FA_cout_1727;
      REGS_829<=FA_cout_1728;
      REGS_830<=FA_cout_1729;
      REGS_831<=FA_cout_1730;
      REGS_832<=FA_cout_1731;
      REGS_833<=FA_cout_1732;
      REGS_834<=FA_cout_1733;
      REGS_835<=FA_cout_1734;
      REGS_836<=FA_cout_1735;
      REGS_837<=FA_cout_1736;
      REGS_838<=FA_cout_1737;
      REGS_839<=FA_cout_1738;
      REGS_840<=FA_cout_1739;
      REGS_841<=FA_cout_1740;
      REGS_842<=FA_cout_1741;
      REGS_843<=FA_cout_1742;
      REGS_844<=FA_cout_1743;
      REGS_845<=FA_cout_1744;
      REGS_846<=FA_cout_1745;
      REGS_847<=FA_cout_1746;
      REGS_848<=FA_cout_1747;
      REGS_849<=FA_cout_1748;
      REGS_850<=FA_cout_1749;
      REGS_851<=FA_cout_1750;
      REGS_852<=FA_cout_1751;
      REGS_853<=FA_out_1752;
      REGS_854<=FA_cout_1752;
      REGS_855<=FA_out_1753;
      REGS_856<=FA_cout_1753;
      REGS_857<=FA_out_1754;
      REGS_858<=FA_cout_1754;
      REGS_859<=FA_out_1755;
      REGS_860<=FA_cout_1755;
      REGS_861<=FA_out_1756;
      REGS_862<=FA_cout_1756;
      REGS_863<=FA_out_1757;
      REGS_864<=FA_cout_1757;
      REGS_865<=FA_out_1716;
      REGS_866<=FA_out_1717;
      REGS_867<=FA_out_1718;
      REGS_868<=FA_out_1719;
      REGS_869<=FA_out_1720;
      REGS_870<=FA_out_1721;
      REGS_871<=FA_out_1722;
      REGS_872<=FA_out_1723;
      REGS_873<=FA_out_1724;
      REGS_874<=FA_out_1725;
      REGS_875<=FA_out_1726;
      REGS_876<=FA_out_1727;
      REGS_877<=FA_out_1728;
      REGS_878<=FA_out_1729;
      REGS_879<=FA_out_1730;
      REGS_880<=FA_out_1731;
      REGS_881<=FA_out_1732;
      REGS_882<=FA_out_1733;
      REGS_883<=FA_out_1734;
      REGS_884<=FA_out_1735;
      REGS_885<=FA_out_1736;
      REGS_886<=FA_out_1737;
      REGS_887<=FA_out_1738;
      REGS_888<=FA_out_1739;
      REGS_889<=FA_out_1740;
      REGS_890<=FA_out_1741;
      REGS_891<=FA_out_1742;
      REGS_892<=FA_out_1743;
      REGS_893<=FA_out_1744;
      REGS_894<=FA_out_1745;
      REGS_895<=FA_out_1746;
      REGS_896<=FA_out_1747;
      REGS_897<=FA_out_1748;
      REGS_898<=FA_out_1749;
      REGS_899<=FA_out_1750;
      REGS_900<=FA_out_1751;
      REGS_901<=FA_out_1758;
      REGS_902<=FA_cout_1758;
      REGS_903<=FA_out_1759;
      REGS_904<=FA_cout_1759;
      REGS_905<=FA_out_1760;
      REGS_906<=FA_cout_1760;
      REGS_907<=FA_out_1761;
      REGS_908<=FA_cout_1761;
      REGS_909<=FA_out_1762;
      REGS_910<=FA_cout_1762;
      REGS_911<=FA_out_1763;
      REGS_912<=FA_cout_1763;
      REGS_913<=FA_out_1764;
      REGS_914<=FA_cout_1764;
      REGS_915<=FA_out_1765;
      REGS_916<=FA_cout_1765;
      REGS_917<=FA_out_1766;
      REGS_918<=FA_cout_1766;
      REGS_919<=FA_out_1767;
      REGS_920<=FA_cout_1767;
      REGS_921<=FA_out_1768;
      REGS_922<=FA_cout_1768;
      REGS_923<=FA_out_1769;
      REGS_924<=FA_cout_1769;
      REGS_925<=FA_out_1770;
      REGS_926<=FA_cout_1770;
      REGS_927<=FA_out_1771;
      REGS_928<=FA_cout_1771;
      REGS_929<=FA_out_1772;
      REGS_930<=FA_cout_1772;
      REGS_931<=FA_out_1773;
      REGS_932<=FA_cout_1773;
      REGS_933<=FA_out_1774;
      REGS_934<=FA_cout_1774;
      REGS_935<=FA_out_1775;
      REGS_936<=FA_cout_1775;
      REGS_937<=FA_out_1776;
      REGS_938<=FA_cout_1776;
      REGS_939<=FA_out_1777;
      REGS_940<=FA_cout_1777;
      REGS_941<=HA_out_52;
      REGS_942<=HA_cout_52;
      REGS_943<=HA_cout_53;
      REGS_944<=HA_cout_54;
      REGS_945<=FA_cout_1778;
      REGS_946<=FA_cout_1779;
      REGS_947<=FA_cout_1780;
      REGS_948<=FA_cout_1781;
      REGS_949<=FA_cout_1782;
      REGS_950<=FA_cout_1783;
      REGS_951<=FA_cout_1784;
      REGS_952<=FA_cout_1785;
      REGS_953<=FA_cout_1786;
      REGS_954<=FA_cout_1787;
      REGS_955<=FA_cout_1788;
      REGS_956<=FA_cout_1789;
      REGS_957<=FA_cout_1790;
      REGS_958<=FA_cout_1791;
      REGS_959<=FA_cout_1792;
      REGS_960<=FA_cout_1793;
      REGS_961<=FA_cout_1794;
      REGS_962<=FA_cout_1795;
      REGS_963<=FA_cout_1796;
      REGS_964<=FA_cout_1797;
      REGS_965<=FA_cout_1798;
      REGS_966<=FA_cout_1799;
      REGS_967<=FA_cout_1800;
      REGS_968<=FA_cout_1801;
      REGS_969<=FA_cout_1802;
      REGS_970<=FA_cout_1803;
      REGS_971<=FA_cout_1804;
      REGS_972<=FA_cout_1805;
      REGS_973<=FA_cout_1806;
      REGS_974<=FA_cout_1807;
      REGS_975<=FA_out_1808;
      REGS_976<=FA_cout_1808;
      REGS_977<=FA_out_1809;
      REGS_978<=FA_cout_1809;
      REGS_979<=FA_out_1810;
      REGS_980<=FA_cout_1810;
      REGS_981<=FA_out_1811;
      REGS_982<=FA_cout_1811;
      REGS_983<=FA_out_1812;
      REGS_984<=FA_cout_1812;
      REGS_985<=FA_out_1813;
      REGS_986<=FA_cout_1813;
      REGS_987<=FA_out_1814;
      REGS_988<=FA_cout_1814;
      REGS_989<=HA_out_53;
      REGS_990<=HA_out_54;
      REGS_991<=FA_out_1778;
      REGS_992<=FA_out_1779;
      REGS_993<=FA_out_1780;
      REGS_994<=FA_out_1781;
      REGS_995<=FA_out_1782;
      REGS_996<=FA_out_1783;
      REGS_997<=FA_out_1784;
      REGS_998<=FA_out_1785;
      REGS_999<=FA_out_1786;
      REGS_1000<=FA_out_1787;
      REGS_1001<=FA_out_1788;
      REGS_1002<=FA_out_1789;
      REGS_1003<=FA_out_1790;
      REGS_1004<=FA_out_1791;
      REGS_1005<=FA_out_1792;
      REGS_1006<=FA_out_1793;
      REGS_1007<=FA_out_1794;
      REGS_1008<=FA_out_1795;
      REGS_1009<=FA_out_1796;
      REGS_1010<=FA_out_1797;
      REGS_1011<=FA_out_1798;
      REGS_1012<=FA_out_1799;
      REGS_1013<=FA_out_1800;
      REGS_1014<=FA_out_1801;
      REGS_1015<=FA_out_1802;
      REGS_1016<=FA_out_1803;
      REGS_1017<=FA_out_1804;
      REGS_1018<=FA_out_1805;
      REGS_1019<=FA_out_1806;
      REGS_1020<=FA_out_1807;
      REGS_1021<=FA_out_1815;
      REGS_1022<=FA_cout_1815;
      REGS_1023<=FA_out_1816;
      REGS_1024<=FA_cout_1816;
      REGS_1025<=FA_out_1817;
      REGS_1026<=FA_cout_1817;
      REGS_1027<=FA_out_1818;
      REGS_1028<=FA_cout_1818;
      REGS_1029<=FA_out_1819;
      REGS_1030<=FA_cout_1819;
      REGS_1031<=FA_out_1820;
      REGS_1032<=FA_cout_1820;
      REGS_1033<=FA_out_1821;
      REGS_1034<=FA_cout_1821;
      REGS_1035<=FA_out_1822;
      REGS_1036<=FA_cout_1822;
      REGS_1037<=FA_out_1823;
      REGS_1038<=FA_cout_1823;
      REGS_1039<=FA_out_1824;
      REGS_1040<=FA_cout_1824;
      REGS_1041<=FA_out_1825;
      REGS_1042<=FA_cout_1825;
      REGS_1043<=FA_out_1826;
      REGS_1044<=FA_cout_1826;
      REGS_1045<=FA_out_1827;
      REGS_1046<=FA_cout_1827;
      REGS_1047<=FA_out_1828;
      REGS_1048<=FA_cout_1828;
      REGS_1049<=FA_out_1829;
      REGS_1050<=FA_cout_1829;
      REGS_1051<=FA_out_1830;
      REGS_1052<=FA_cout_1830;
      REGS_1053<=FA_out_1831;
      REGS_1054<=FA_cout_1831;
      REGS_1055<=FA_out_1832;
      REGS_1056<=FA_cout_1832;
      REGS_1057<=FA_out_1833;
      REGS_1058<=FA_cout_1833;
      REGS_1059<=FA_out_1834;
      REGS_1060<=FA_cout_1834;
      REGS_1061<=FA_out_1835;
      REGS_1062<=FA_cout_1835;
      REGS_1063<=FA_out_1836;
      REGS_1064<=FA_cout_1836;
      REGS_1065<=FA_out_1837;
      REGS_1066<=FA_cout_1837;
      REGS_1067<=FA_out_1838;
      REGS_1068<=FA_cout_1838;
      REGS_1069<=FA_out_1839;
      REGS_1070<=FA_cout_1839;
      REGS_1071<=FA_out_1840;
      REGS_1072<=FA_cout_1840;
      REGS_1073<=FA_out_1841;
      REGS_1074<=FA_cout_1841;
      REGS_1075<=FA_out_1842;
      REGS_1076<=FA_cout_1842;
      REGS_1077<=FA_out_1843;
      REGS_1078<=FA_cout_1843;
      REGS_1079<=FA_out_1844;
      REGS_1080<=FA_cout_1844;
      REGS_1081<=FA_out_1845;
      REGS_1082<=FA_cout_1845;
      REGS_1083<=FA_out_1846;
      REGS_1084<=FA_cout_1846;
      REGS_1085<=inp_36[0];
      REGS_1086<=HA_out_12;
      REGS_1087<=HA_out_55;
      REGS_1088<=HA_cout_55;
      REGS_1089<=FA_cout_1847;
      REGS_1090<=FA_cout_1848;
      REGS_1091<=FA_cout_1849;
      REGS_1092<=FA_cout_1850;
      REGS_1093<=FA_cout_1851;
      REGS_1094<=FA_cout_1852;
      REGS_1095<=FA_cout_1853;
      REGS_1096<=FA_cout_1854;
      REGS_1097<=FA_cout_1855;
      REGS_1098<=FA_cout_1856;
      REGS_1099<=FA_cout_1857;
      REGS_1100<=FA_cout_1858;
      REGS_1101<=FA_cout_1859;
      REGS_1102<=FA_cout_1860;
      REGS_1103<=FA_cout_1861;
      REGS_1104<=FA_cout_1862;
      REGS_1105<=FA_cout_1863;
      REGS_1106<=FA_cout_1864;
      REGS_1107<=FA_cout_1865;
      REGS_1108<=FA_cout_1866;
      REGS_1109<=FA_cout_1867;
      REGS_1110<=FA_cout_1868;
      REGS_1111<=FA_cout_1869;
      REGS_1112<=FA_cout_1870;
      REGS_1113<=FA_cout_1871;
      REGS_1114<=FA_cout_1872;
      REGS_1115<=FA_cout_1873;
      REGS_1116<=FA_out_1874;
      REGS_1117<=FA_cout_1874;
      REGS_1118<=FA_out_1875;
      REGS_1119<=FA_cout_1875;
      REGS_1120<=FA_out_1876;
      REGS_1121<=FA_cout_1876;
      REGS_1122<=FA_out_1877;
      REGS_1123<=FA_cout_1877;
      REGS_1124<=FA_out_1878;
      REGS_1125<=FA_cout_1878;
      REGS_1126<=FA_out_1879;
      REGS_1127<=FA_cout_1879;
      REGS_1128<=FA_out_1880;
      REGS_1129<=FA_cout_1880;
      REGS_1130<=FA_out_1881;
      REGS_1131<=FA_cout_1881;
      REGS_1132<=FA_out_1847;
      REGS_1133<=FA_out_1848;
      REGS_1134<=FA_out_1849;
      REGS_1135<=FA_out_1850;
      REGS_1136<=FA_out_1851;
      REGS_1137<=FA_out_1852;
      REGS_1138<=FA_out_1853;
      REGS_1139<=FA_out_1854;
      REGS_1140<=FA_out_1855;
      REGS_1141<=FA_out_1856;
      REGS_1142<=FA_out_1857;
      REGS_1143<=FA_out_1858;
      REGS_1144<=FA_out_1859;
      REGS_1145<=FA_out_1860;
      REGS_1146<=FA_out_1861;
      REGS_1147<=FA_out_1862;
      REGS_1148<=FA_out_1863;
      REGS_1149<=FA_out_1864;
      REGS_1150<=FA_out_1865;
      REGS_1151<=FA_out_1866;
      REGS_1152<=FA_out_1867;
      REGS_1153<=FA_out_1868;
      REGS_1154<=FA_out_1869;
      REGS_1155<=FA_out_1870;
      REGS_1156<=FA_out_1871;
      REGS_1157<=FA_out_1872;
      REGS_1158<=FA_out_1873;
      REGS_1159<=FA_out_1882;
      REGS_1160<=FA_cout_1882;
      REGS_1161<=FA_out_1883;
      REGS_1162<=FA_cout_1883;
      REGS_1163<=FA_out_1884;
      REGS_1164<=FA_cout_1884;
      REGS_1165<=FA_out_1885;
      REGS_1166<=FA_cout_1885;
      REGS_1167<=FA_out_1886;
      REGS_1168<=FA_cout_1886;
      REGS_1169<=FA_out_1887;
      REGS_1170<=FA_cout_1887;
      REGS_1171<=FA_out_1888;
      REGS_1172<=FA_cout_1888;
      REGS_1173<=FA_out_1889;
      REGS_1174<=FA_cout_1889;
      REGS_1175<=FA_out_1890;
      REGS_1176<=FA_cout_1890;
      REGS_1177<=FA_out_1891;
      REGS_1178<=FA_cout_1891;
      REGS_1179<=FA_out_1892;
      REGS_1180<=FA_cout_1892;
      REGS_1181<=FA_out_1893;
      REGS_1182<=FA_cout_1893;
      REGS_1183<=FA_out_1894;
      REGS_1184<=FA_cout_1894;
      REGS_1185<=FA_out_1895;
      REGS_1186<=FA_cout_1895;
      REGS_1187<=FA_out_1896;
      REGS_1188<=FA_cout_1896;
      REGS_1189<=FA_out_1897;
      REGS_1190<=FA_cout_1897;
      REGS_1191<=FA_out_1898;
      REGS_1192<=FA_cout_1898;
      REGS_1193<=FA_out_1899;
      REGS_1194<=FA_cout_1899;
      REGS_1195<=FA_out_1900;
      REGS_1196<=FA_cout_1900;
      REGS_1197<=FA_out_1901;
      REGS_1198<=FA_cout_1901;
      REGS_1199<=FA_out_1902;
      REGS_1200<=FA_cout_1902;
      REGS_1201<=FA_out_1903;
      REGS_1202<=FA_cout_1903;
      REGS_1203<=FA_out_1904;
      REGS_1204<=FA_cout_1904;
      REGS_1205<=FA_out_1905;
      REGS_1206<=FA_cout_1905;
      REGS_1207<=FA_out_1906;
      REGS_1208<=FA_cout_1906;
      REGS_1209<=FA_out_1907;
      REGS_1210<=FA_cout_1907;
      REGS_1211<=FA_out_832;
      REGS_1212<=HA_out_56;
      REGS_1213<=HA_cout_56;
      REGS_1214<=HA_cout_57;
      REGS_1215<=FA_cout_1908;
      REGS_1216<=FA_cout_1909;
      REGS_1217<=FA_cout_1910;
      REGS_1218<=FA_cout_1911;
      REGS_1219<=FA_cout_1912;
      REGS_1220<=FA_cout_1913;
      REGS_1221<=FA_cout_1914;
      REGS_1222<=FA_cout_1915;
      REGS_1223<=FA_cout_1916;
      REGS_1224<=FA_cout_1917;
      REGS_1225<=FA_cout_1918;
      REGS_1226<=FA_cout_1919;
      REGS_1227<=FA_cout_1920;
      REGS_1228<=FA_cout_1921;
      REGS_1229<=FA_cout_1922;
      REGS_1230<=FA_cout_1923;
      REGS_1231<=FA_cout_1924;
      REGS_1232<=FA_cout_1925;
      REGS_1233<=FA_cout_1926;
      REGS_1234<=FA_cout_1927;
      REGS_1235<=FA_cout_1928;
      REGS_1236<=FA_out_1929;
      REGS_1237<=FA_cout_1929;
      REGS_1238<=FA_out_1930;
      REGS_1239<=FA_cout_1930;
      REGS_1240<=FA_out_1931;
      REGS_1241<=FA_cout_1931;
      REGS_1242<=FA_out_1932;
      REGS_1243<=FA_cout_1932;
      REGS_1244<=FA_out_1933;
      REGS_1245<=FA_cout_1933;
      REGS_1246<=FA_out_1934;
      REGS_1247<=FA_cout_1934;
      REGS_1248<=FA_out_1935;
      REGS_1249<=FA_cout_1935;
      REGS_1250<=FA_out_1936;
      REGS_1251<=FA_cout_1936;
      REGS_1252<=FA_out_1937;
      REGS_1253<=FA_cout_1937;
      REGS_1254<=HA_out_57;
      REGS_1255<=FA_out_1908;
      REGS_1256<=FA_out_1909;
      REGS_1257<=FA_out_1910;
      REGS_1258<=FA_out_1911;
      REGS_1259<=FA_out_1912;
      REGS_1260<=FA_out_1913;
      REGS_1261<=FA_out_1914;
      REGS_1262<=FA_out_1915;
      REGS_1263<=FA_out_1916;
      REGS_1264<=FA_out_1917;
      REGS_1265<=FA_out_1918;
      REGS_1266<=FA_out_1919;
      REGS_1267<=FA_out_1920;
      REGS_1268<=FA_out_1921;
      REGS_1269<=FA_out_1922;
      REGS_1270<=FA_out_1923;
      REGS_1271<=FA_out_1924;
      REGS_1272<=FA_out_1925;
      REGS_1273<=FA_out_1926;
      REGS_1274<=FA_out_1927;
      REGS_1275<=FA_out_1928;
      REGS_1276<=FA_out_1938;
      REGS_1277<=FA_cout_1938;
      REGS_1278<=FA_out_1939;
      REGS_1279<=FA_cout_1939;
      REGS_1280<=FA_out_1940;
      REGS_1281<=FA_cout_1940;
      REGS_1282<=FA_out_1941;
      REGS_1283<=FA_cout_1941;
      REGS_1284<=FA_out_1942;
      REGS_1285<=FA_cout_1942;
      REGS_1286<=FA_out_1943;
      REGS_1287<=FA_cout_1943;
      REGS_1288<=FA_out_1944;
      REGS_1289<=FA_cout_1944;
      REGS_1290<=FA_out_1945;
      REGS_1291<=FA_cout_1945;
      REGS_1292<=FA_out_1946;
      REGS_1293<=FA_cout_1946;
      REGS_1294<=FA_out_1947;
      REGS_1295<=FA_cout_1947;
      REGS_1296<=FA_out_1948;
      REGS_1297<=FA_cout_1948;
      REGS_1298<=FA_out_1949;
      REGS_1299<=FA_cout_1949;
      REGS_1300<=FA_out_1950;
      REGS_1301<=FA_cout_1950;
      REGS_1302<=FA_out_1951;
      REGS_1303<=FA_cout_1951;
      REGS_1304<=FA_out_1952;
      REGS_1305<=FA_cout_1952;
      REGS_1306<=FA_out_1953;
      REGS_1307<=FA_cout_1953;
      REGS_1308<=FA_out_1954;
      REGS_1309<=FA_cout_1954;
      REGS_1310<=FA_out_1955;
      REGS_1311<=FA_cout_1955;
      REGS_1312<=FA_out_1956;
      REGS_1313<=FA_cout_1956;
      REGS_1314<=FA_out_1957;
      REGS_1315<=FA_cout_1957;
      REGS_1316<=FA_out_1958;
      REGS_1317<=FA_cout_1958;
      REGS_1318<=FA_out_1959;
      REGS_1319<=FA_cout_1959;
      REGS_1320<=FA_out_1960;
      REGS_1321<=FA_cout_1960;
      REGS_1322<=FA_out_1961;
      REGS_1323<=FA_cout_1961;
      REGS_1324<=FA_out_1962;
      REGS_1325<=FA_cout_1962;
      REGS_1326<=FA_out_1963;
      REGS_1327<=FA_cout_1963;
      REGS_1328<=FA_out_1964;
      REGS_1329<=FA_cout_1964;
      REGS_1330<=FA_out_1965;
      REGS_1331<=FA_cout_1965;
      REGS_1332<=FA_out_1966;
      REGS_1333<=FA_cout_1966;
      REGS_1334<=FA_out_1967;
      REGS_1335<=FA_cout_1967;
      REGS_1336<=FA_out_1968;
      REGS_1337<=FA_cout_1968;
      REGS_1338<=FA_out_1969;
      REGS_1339<=FA_cout_1969;
      REGS_1340<=FA_out_1970;
      REGS_1341<=FA_cout_1970;
      REGS_1342<=FA_out_1971;
      REGS_1343<=FA_cout_1971;
      REGS_1344<=FA_out_1972;
      REGS_1345<=FA_cout_1972;
      REGS_1346<=FA_out_1973;
      REGS_1347<=FA_cout_1973;
      REGS_1348<=FA_out_1974;
      REGS_1349<=FA_cout_1974;
      REGS_1350<=FA_out_1975;
      REGS_1351<=FA_cout_1975;
      REGS_1352<=FA_out_1976;
      REGS_1353<=FA_cout_1976;
      REGS_1354<=FA_out_1977;
      REGS_1355<=FA_cout_1977;
      REGS_1356<=inp_45[0];
      REGS_1357<=HA_out_15;
      REGS_1358<=HA_out_58;
      REGS_1359<=HA_cout_58;
      REGS_1360<=FA_cout_1978;
      REGS_1361<=FA_cout_1979;
      REGS_1362<=FA_cout_1980;
      REGS_1363<=FA_cout_1981;
      REGS_1364<=FA_cout_1982;
      REGS_1365<=FA_cout_1983;
      REGS_1366<=FA_cout_1984;
      REGS_1367<=FA_cout_1985;
      REGS_1368<=FA_cout_1986;
      REGS_1369<=FA_cout_1987;
      REGS_1370<=FA_cout_1988;
      REGS_1371<=FA_cout_1989;
      REGS_1372<=FA_cout_1990;
      REGS_1373<=FA_cout_1991;
      REGS_1374<=FA_cout_1992;
      REGS_1375<=FA_cout_1993;
      REGS_1376<=FA_cout_1994;
      REGS_1377<=FA_cout_1995;
      REGS_1378<=FA_out_1996;
      REGS_1379<=FA_cout_1996;
      REGS_1380<=FA_out_1997;
      REGS_1381<=FA_cout_1997;
      REGS_1382<=FA_out_1998;
      REGS_1383<=FA_cout_1998;
      REGS_1384<=FA_out_1999;
      REGS_1385<=FA_cout_1999;
      REGS_1386<=FA_out_2000;
      REGS_1387<=FA_cout_2000;
      REGS_1388<=FA_out_2001;
      REGS_1389<=FA_cout_2001;
      REGS_1390<=FA_out_2002;
      REGS_1391<=FA_cout_2002;
      REGS_1392<=FA_out_2003;
      REGS_1393<=FA_cout_2003;
      REGS_1394<=FA_out_2004;
      REGS_1395<=FA_cout_2004;
      REGS_1396<=FA_out_2005;
      REGS_1397<=FA_cout_2005;
      REGS_1398<=FA_out_1978;
      REGS_1399<=FA_out_1979;
      REGS_1400<=FA_out_1980;
      REGS_1401<=FA_out_1981;
      REGS_1402<=FA_out_1982;
      REGS_1403<=FA_out_1983;
      REGS_1404<=FA_out_1984;
      REGS_1405<=FA_out_1985;
      REGS_1406<=FA_out_1986;
      REGS_1407<=FA_out_1987;
      REGS_1408<=FA_out_1988;
      REGS_1409<=FA_out_1989;
      REGS_1410<=FA_out_1990;
      REGS_1411<=FA_out_1991;
      REGS_1412<=FA_out_1992;
      REGS_1413<=FA_out_1993;
      REGS_1414<=FA_out_1994;
      REGS_1415<=FA_out_1995;
      REGS_1416<=FA_out_2006;
      REGS_1417<=FA_cout_2006;
      REGS_1418<=FA_out_2007;
      REGS_1419<=FA_cout_2007;
      REGS_1420<=FA_out_2008;
      REGS_1421<=FA_cout_2008;
      REGS_1422<=FA_out_2009;
      REGS_1423<=FA_cout_2009;
      REGS_1424<=FA_out_2010;
      REGS_1425<=FA_cout_2010;
      REGS_1426<=FA_out_2011;
      REGS_1427<=FA_cout_2011;
      REGS_1428<=FA_out_2012;
      REGS_1429<=FA_cout_2012;
      REGS_1430<=FA_out_2013;
      REGS_1431<=FA_cout_2013;
      REGS_1432<=FA_out_2014;
      REGS_1433<=FA_cout_2014;
      REGS_1434<=FA_out_2015;
      REGS_1435<=FA_cout_2015;
      REGS_1436<=FA_out_2016;
      REGS_1437<=FA_cout_2016;
      REGS_1438<=FA_out_2017;
      REGS_1439<=FA_cout_2017;
      REGS_1440<=FA_out_2018;
      REGS_1441<=FA_cout_2018;
      REGS_1442<=FA_out_2019;
      REGS_1443<=FA_cout_2019;
      REGS_1444<=FA_out_2020;
      REGS_1445<=FA_cout_2020;
      REGS_1446<=FA_out_2021;
      REGS_1447<=FA_cout_2021;
      REGS_1448<=FA_out_2022;
      REGS_1449<=FA_cout_2022;
      REGS_1450<=FA_out_2023;
      REGS_1451<=FA_cout_2023;
      REGS_1452<=FA_out_2024;
      REGS_1453<=FA_cout_2024;
      REGS_1454<=FA_out_2025;
      REGS_1455<=FA_cout_2025;
      REGS_1456<=FA_out_2026;
      REGS_1457<=FA_cout_2026;
      REGS_1458<=FA_out_2027;
      REGS_1459<=FA_cout_2027;
      REGS_1460<=FA_out_2028;
      REGS_1461<=FA_cout_2028;
      REGS_1462<=FA_out_2029;
      REGS_1463<=FA_cout_2029;
      REGS_1464<=FA_out_2030;
      REGS_1465<=FA_cout_2030;
      REGS_1466<=FA_out_2031;
      REGS_1467<=FA_cout_2031;
      REGS_1468<=FA_out_2032;
      REGS_1469<=FA_cout_2032;
      REGS_1470<=FA_out_2033;
      REGS_1471<=FA_cout_2033;
      REGS_1472<=FA_out_2034;
      REGS_1473<=FA_cout_2034;
      REGS_1474<=FA_out_2035;
      REGS_1475<=FA_cout_2035;
      REGS_1476<=FA_out_2036;
      REGS_1477<=FA_cout_2036;
      REGS_1478<=FA_out_2037;
      REGS_1479<=FA_cout_2037;
      REGS_1480<=FA_out_1024;
      REGS_1481<=HA_out_59;
      REGS_1482<=HA_cout_59;
      REGS_1483<=HA_cout_60;
      REGS_1484<=FA_cout_2038;
      REGS_1485<=FA_cout_2039;
      REGS_1486<=FA_cout_2040;
      REGS_1487<=FA_cout_2041;
      REGS_1488<=FA_cout_2042;
      REGS_1489<=FA_cout_2043;
      REGS_1490<=FA_cout_2044;
      REGS_1491<=FA_cout_2045;
      REGS_1492<=FA_cout_2046;
      REGS_1493<=FA_cout_2047;
      REGS_1494<=FA_cout_2048;
      REGS_1495<=FA_cout_2049;
      REGS_1496<=FA_out_2050;
      REGS_1497<=FA_cout_2050;
      REGS_1498<=FA_out_2051;
      REGS_1499<=FA_cout_2051;
      REGS_1500<=FA_out_2052;
      REGS_1501<=FA_cout_2052;
      REGS_1502<=FA_out_2053;
      REGS_1503<=FA_cout_2053;
      REGS_1504<=FA_out_2054;
      REGS_1505<=FA_cout_2054;
      REGS_1506<=FA_out_2055;
      REGS_1507<=FA_cout_2055;
      REGS_1508<=FA_out_2056;
      REGS_1509<=FA_cout_2056;
      REGS_1510<=FA_out_2057;
      REGS_1511<=FA_cout_2057;
      REGS_1512<=FA_out_2058;
      REGS_1513<=FA_cout_2058;
      REGS_1514<=FA_out_2059;
      REGS_1515<=FA_cout_2059;
      REGS_1516<=FA_out_2060;
      REGS_1517<=FA_cout_2060;
      REGS_1518<=HA_out_60;
      REGS_1519<=FA_out_2038;
      REGS_1520<=FA_out_2039;
      REGS_1521<=FA_out_2040;
      REGS_1522<=FA_out_2041;
      REGS_1523<=FA_out_2042;
      REGS_1524<=FA_out_2043;
      REGS_1525<=FA_out_2044;
      REGS_1526<=FA_out_2045;
      REGS_1527<=FA_out_2046;
      REGS_1528<=FA_out_2047;
      REGS_1529<=FA_out_2048;
      REGS_1530<=FA_out_2049;
      REGS_1531<=FA_out_2061;
      REGS_1532<=FA_cout_2061;
      REGS_1533<=FA_out_2062;
      REGS_1534<=FA_cout_2062;
      REGS_1535<=FA_out_2063;
      REGS_1536<=FA_cout_2063;
      REGS_1537<=FA_out_2064;
      REGS_1538<=FA_cout_2064;
      REGS_1539<=FA_out_2065;
      REGS_1540<=FA_cout_2065;
      REGS_1541<=FA_out_2066;
      REGS_1542<=FA_cout_2066;
      REGS_1543<=FA_out_2067;
      REGS_1544<=FA_cout_2067;
      REGS_1545<=FA_out_2068;
      REGS_1546<=FA_cout_2068;
      REGS_1547<=FA_out_2069;
      REGS_1548<=FA_cout_2069;
      REGS_1549<=FA_out_2070;
      REGS_1550<=FA_cout_2070;
      REGS_1551<=FA_out_2071;
      REGS_1552<=FA_cout_2071;
      REGS_1553<=FA_out_2072;
      REGS_1554<=FA_cout_2072;
      REGS_1555<=FA_out_2073;
      REGS_1556<=FA_cout_2073;
      REGS_1557<=FA_out_2074;
      REGS_1558<=FA_cout_2074;
      REGS_1559<=FA_out_2075;
      REGS_1560<=FA_cout_2075;
      REGS_1561<=FA_out_2076;
      REGS_1562<=FA_cout_2076;
      REGS_1563<=FA_out_2077;
      REGS_1564<=FA_cout_2077;
      REGS_1565<=FA_out_2078;
      REGS_1566<=FA_cout_2078;
      REGS_1567<=FA_out_2079;
      REGS_1568<=FA_cout_2079;
      REGS_1569<=FA_out_2080;
      REGS_1570<=FA_cout_2080;
      REGS_1571<=FA_out_2081;
      REGS_1572<=FA_cout_2081;
      REGS_1573<=FA_out_2082;
      REGS_1574<=FA_cout_2082;
      REGS_1575<=FA_out_2083;
      REGS_1576<=FA_cout_2083;
      REGS_1577<=FA_out_2084;
      REGS_1578<=FA_cout_2084;
      REGS_1579<=FA_out_2085;
      REGS_1580<=FA_cout_2085;
      REGS_1581<=FA_out_2086;
      REGS_1582<=FA_cout_2086;
      REGS_1583<=FA_out_2087;
      REGS_1584<=FA_cout_2087;
      REGS_1585<=FA_out_2088;
      REGS_1586<=FA_cout_2088;
      REGS_1587<=FA_out_2089;
      REGS_1588<=FA_cout_2089;
      REGS_1589<=FA_out_2090;
      REGS_1590<=FA_cout_2090;
      REGS_1591<=FA_out_2091;
      REGS_1592<=FA_cout_2091;
      REGS_1593<=FA_out_2092;
      REGS_1594<=FA_cout_2092;
      REGS_1595<=FA_out_2093;
      REGS_1596<=FA_cout_2093;
      REGS_1597<=FA_out_2094;
      REGS_1598<=FA_cout_2094;
      REGS_1599<=FA_out_2095;
      REGS_1600<=FA_cout_2095;
      REGS_1601<=FA_out_2096;
      REGS_1602<=FA_cout_2096;
      REGS_1603<=FA_out_2097;
      REGS_1604<=FA_cout_2097;
      REGS_1605<=FA_out_2098;
      REGS_1606<=FA_cout_2098;
      REGS_1607<=FA_out_2099;
      REGS_1608<=FA_cout_2099;
      REGS_1609<=FA_out_2100;
      REGS_1610<=FA_cout_2100;
      REGS_1611<=FA_out_2101;
      REGS_1612<=FA_cout_2101;
      REGS_1613<=FA_out_2102;
      REGS_1614<=FA_cout_2102;
      REGS_1615<=FA_out_2103;
      REGS_1616<=FA_cout_2103;
      REGS_1617<=FA_out_2104;
      REGS_1618<=FA_cout_2104;
      REGS_1619<=FA_out_2105;
      REGS_1620<=FA_cout_2105;
      REGS_1621<=FA_out_2106;
      REGS_1622<=FA_cout_2106;
      REGS_1623<=FA_out_2107;
      REGS_1624<=FA_cout_2107;
      REGS_1625<=FA_out_2108;
      REGS_1626<=FA_cout_2108;
      REGS_1627<=inp_54[0];
      REGS_1628<=HA_out_18;
      REGS_1629<=HA_out_61;
      REGS_1630<=HA_cout_61;
      REGS_1631<=FA_cout_2109;
      REGS_1632<=FA_cout_2110;
      REGS_1633<=FA_cout_2111;
      REGS_1634<=FA_cout_2112;
      REGS_1635<=FA_cout_2113;
      REGS_1636<=FA_cout_2114;
      REGS_1637<=FA_cout_2115;
      REGS_1638<=FA_cout_2116;
      REGS_1639<=FA_cout_2117;
      REGS_1640<=FA_out_2118;
      REGS_1641<=FA_cout_2118;
      REGS_1642<=FA_out_2119;
      REGS_1643<=FA_cout_2119;
      REGS_1644<=FA_out_2120;
      REGS_1645<=FA_cout_2120;
      REGS_1646<=FA_out_2121;
      REGS_1647<=FA_cout_2121;
      REGS_1648<=FA_out_2122;
      REGS_1649<=FA_cout_2122;
      REGS_1650<=FA_out_2123;
      REGS_1651<=FA_cout_2123;
      REGS_1652<=FA_out_2124;
      REGS_1653<=FA_cout_2124;
      REGS_1654<=FA_out_2125;
      REGS_1655<=FA_cout_2125;
      REGS_1656<=FA_out_2126;
      REGS_1657<=FA_cout_2126;
      REGS_1658<=FA_out_2127;
      REGS_1659<=FA_cout_2127;
      REGS_1660<=FA_out_2128;
      REGS_1661<=FA_cout_2128;
      REGS_1662<=FA_out_2129;
      REGS_1663<=FA_cout_2129;
      REGS_1664<=FA_out_2109;
      REGS_1665<=FA_out_2110;
      REGS_1666<=FA_out_2111;
      REGS_1667<=FA_out_2112;
      REGS_1668<=FA_out_2113;
      REGS_1669<=FA_out_2114;
      REGS_1670<=FA_out_2115;
      REGS_1671<=FA_out_2116;
      REGS_1672<=FA_out_2117;
      REGS_1673<=FA_out_2130;
      REGS_1674<=FA_cout_2130;
      REGS_1675<=FA_out_2131;
      REGS_1676<=FA_cout_2131;
      REGS_1677<=FA_out_2132;
      REGS_1678<=FA_cout_2132;
      REGS_1679<=FA_out_2133;
      REGS_1680<=FA_cout_2133;
      REGS_1681<=FA_out_2134;
      REGS_1682<=FA_cout_2134;
      REGS_1683<=FA_out_2135;
      REGS_1684<=FA_cout_2135;
      REGS_1685<=FA_out_2136;
      REGS_1686<=FA_cout_2136;
      REGS_1687<=FA_out_2137;
      REGS_1688<=FA_cout_2137;
      REGS_1689<=FA_out_2138;
      REGS_1690<=FA_cout_2138;
      REGS_1691<=FA_out_2139;
      REGS_1692<=FA_cout_2139;
      REGS_1693<=FA_out_2140;
      REGS_1694<=FA_cout_2140;
      REGS_1695<=FA_out_2141;
      REGS_1696<=FA_cout_2141;
      REGS_1697<=FA_out_2142;
      REGS_1698<=FA_cout_2142;
      REGS_1699<=FA_out_2143;
      REGS_1700<=FA_cout_2143;
      REGS_1701<=FA_out_2144;
      REGS_1702<=FA_cout_2144;
      REGS_1703<=FA_out_2145;
      REGS_1704<=FA_cout_2145;
      REGS_1705<=FA_out_2146;
      REGS_1706<=FA_cout_2146;
      REGS_1707<=FA_out_2147;
      REGS_1708<=FA_cout_2147;
      REGS_1709<=FA_out_2148;
      REGS_1710<=FA_cout_2148;
      REGS_1711<=FA_out_2149;
      REGS_1712<=FA_cout_2149;
      REGS_1713<=FA_out_2150;
      REGS_1714<=FA_cout_2150;
      REGS_1715<=FA_out_2151;
      REGS_1716<=FA_cout_2151;
      REGS_1717<=FA_out_2152;
      REGS_1718<=FA_cout_2152;
      REGS_1719<=FA_out_2153;
      REGS_1720<=FA_cout_2153;
      REGS_1721<=FA_out_2154;
      REGS_1722<=FA_cout_2154;
      REGS_1723<=FA_out_2155;
      REGS_1724<=FA_cout_2155;
      REGS_1725<=FA_out_2156;
      REGS_1726<=FA_cout_2156;
      REGS_1727<=FA_out_2157;
      REGS_1728<=FA_cout_2157;
      REGS_1729<=FA_out_2158;
      REGS_1730<=FA_cout_2158;
      REGS_1731<=FA_out_2159;
      REGS_1732<=FA_cout_2159;
      REGS_1733<=FA_out_2160;
      REGS_1734<=FA_cout_2160;
      REGS_1735<=FA_out_2161;
      REGS_1736<=FA_cout_2161;
      REGS_1737<=FA_out_2162;
      REGS_1738<=FA_cout_2162;
      REGS_1739<=FA_out_2163;
      REGS_1740<=FA_cout_2163;
      REGS_1741<=FA_out_2164;
      REGS_1742<=FA_cout_2164;
      REGS_1743<=FA_out_2165;
      REGS_1744<=FA_cout_2165;
      REGS_1745<=FA_out_2166;
      REGS_1746<=FA_cout_2166;
      REGS_1747<=FA_out_2167;
      REGS_1748<=FA_cout_2167;
      REGS_1749<=FA_out_1216;
      REGS_1750<=HA_out_62;
      REGS_1751<=HA_cout_62;
      REGS_1752<=HA_cout_63;
      REGS_1753<=FA_cout_2168;
      REGS_1754<=FA_cout_2169;
      REGS_1755<=FA_cout_2170;
      REGS_1756<=FA_out_2171;
      REGS_1757<=FA_cout_2171;
      REGS_1758<=FA_out_2172;
      REGS_1759<=FA_cout_2172;
      REGS_1760<=FA_out_2173;
      REGS_1761<=FA_cout_2173;
      REGS_1762<=FA_out_2174;
      REGS_1763<=FA_cout_2174;
      REGS_1764<=FA_out_2175;
      REGS_1765<=FA_cout_2175;
      REGS_1766<=FA_out_2176;
      REGS_1767<=FA_cout_2176;
      REGS_1768<=FA_out_2177;
      REGS_1769<=FA_cout_2177;
      REGS_1770<=FA_out_2178;
      REGS_1771<=FA_cout_2178;
      REGS_1772<=FA_out_2179;
      REGS_1773<=FA_cout_2179;
      REGS_1774<=FA_out_2180;
      REGS_1775<=FA_cout_2180;
      REGS_1776<=FA_out_2181;
      REGS_1777<=FA_cout_2181;
      REGS_1778<=FA_out_2182;
      REGS_1779<=FA_cout_2182;
      REGS_1780<=FA_out_2183;
      REGS_1781<=FA_cout_2183;
      REGS_1782<=HA_out_63;
      REGS_1783<=FA_out_2168;
      REGS_1784<=FA_out_2169;
      REGS_1785<=FA_out_2170;
      REGS_1786<=FA_out_2184;
      REGS_1787<=FA_cout_2184;
      REGS_1788<=FA_out_2185;
      REGS_1789<=FA_cout_2185;
      REGS_1790<=FA_out_2186;
      REGS_1791<=FA_cout_2186;
      REGS_1792<=FA_out_2187;
      REGS_1793<=FA_cout_2187;
      REGS_1794<=FA_out_2188;
      REGS_1795<=FA_cout_2188;
      REGS_1796<=FA_out_2189;
      REGS_1797<=FA_cout_2189;
      REGS_1798<=FA_out_2190;
      REGS_1799<=FA_cout_2190;
      REGS_1800<=FA_out_2191;
      REGS_1801<=FA_cout_2191;
      REGS_1802<=FA_out_2192;
      REGS_1803<=FA_cout_2192;
      REGS_1804<=FA_out_2193;
      REGS_1805<=FA_cout_2193;
      REGS_1806<=FA_out_2194;
      REGS_1807<=FA_cout_2194;
      REGS_1808<=FA_out_2195;
      REGS_1809<=FA_cout_2195;
      REGS_1810<=FA_out_2196;
      REGS_1811<=FA_cout_2196;
      REGS_1812<=FA_out_2197;
      REGS_1813<=FA_cout_2197;
      REGS_1814<=FA_out_2198;
      REGS_1815<=FA_cout_2198;
      REGS_1816<=HA_out_64;
      REGS_1817<=HA_cout_64;
      REGS_1818<=FA_out_2199;
      REGS_1819<=FA_cout_2199;
      REGS_1820<=HA_out_65;
      REGS_1821<=HA_cout_65;
      REGS_1822<=FA_out_2200;
      REGS_1823<=FA_cout_2200;
      REGS_1824<=HA_out_66;
      REGS_1825<=HA_cout_66;
      REGS_1826<=FA_out_2201;
      REGS_1827<=FA_cout_2201;
      REGS_1828<=HA_out_67;
      REGS_1829<=HA_cout_67;
      REGS_1830<=FA_out_2202;
      REGS_1831<=FA_cout_2202;
      REGS_1832<=HA_out_68;
      REGS_1833<=HA_cout_68;
      REGS_1834<=FA_out_2203;
      REGS_1835<=FA_cout_2203;
      REGS_1836<=HA_out_69;
      REGS_1837<=HA_cout_69;
      REGS_1838<=FA_out_2204;
      REGS_1839<=FA_cout_2204;
      REGS_1840<=HA_out_70;
      REGS_1841<=HA_cout_70;
      REGS_1842<=FA_out_1303;
      REGS_1843<=HA_out_71;
      REGS_1844<=HA_cout_71;
      REGS_1845<=FA_out_1306;
      REGS_1846<=HA_out_72;
      REGS_1847<=HA_cout_72;
      REGS_1848<=FA_out_1309;
      REGS_1849<=HA_out_73;
      REGS_1850<=HA_cout_73;
      REGS_1851<=FA_out_1312;
      REGS_1852<=HA_out_74;
      REGS_1853<=HA_cout_74;
      REGS_1854<=FA_out_1315;
      REGS_1855<=HA_out_75;
      REGS_1856<=HA_cout_75;
      REGS_1857<=FA_out_1318;
      REGS_1858<=HA_out_76;
      REGS_1859<=HA_cout_76;
      REGS_1860<=FA_out_1321;
      REGS_1861<=HA_out_77;
      REGS_1862<=HA_cout_77;
      REGS_1863<=HA_out_22;
      REGS_1864<=HA_out_78;
      REGS_1865<=HA_cout_78;
      REGS_1866<=HA_out_25;
      REGS_1867<=HA_out_79;
      REGS_1868<=HA_cout_79;
      REGS_1869<=HA_out_28;
      REGS_1870<=HA_out_80;
      REGS_1871<=HA_cout_80;
      REGS_1872<=HA_out_31;
      REGS_1873<=HA_out_81;
      REGS_1874<=HA_cout_81;
      REGS_1875<=HA_out_34;
      REGS_1876<=HA_out_82;
      REGS_1877<=HA_cout_82;
      REGS_1878<=HA_out_37;
      REGS_1879<=HA_out_83;
      REGS_1880<=HA_cout_83;
      REGS_1881<=HA_out_40;
      REGS_1882<=HA_out_84;
      REGS_1883<=HA_cout_84;
      REGS_1884<=inp_63[0];
      REGS_1885<=inp_63[1];
      REGS_1886<=inp_63[6];
      REGS_1887<=inp_63[15];
      REGS_1888<=inp_63[24];
      REGS_1889<=inp_63[33];
      REGS_1890<=inp_63[42];
      REGS_1891<=inp_63[51];
      REGS_1892<=inp_63[60];
      REGS_1893<=REGS_0;
      REGS_1894<=REGS_1;
      REGS_1895<=REGS_2;
      REGS_1896<=HA_out_85;
      REGS_1897<=HA_out_128;
      REGS_1898<=HA_out_171;
      REGS_1899<=HA_out_215;
      REGS_1900<=HA_cout_215;
      REGS_1901<=HA_cout_216;
      REGS_1902<=HA_cout_217;
      REGS_1903<=HA_cout_218;
      REGS_1904<=HA_cout_219;
      REGS_1905<=HA_cout_220;
      REGS_1906<=HA_cout_221;
      REGS_1907<=HA_cout_222;
      REGS_1908<=HA_cout_223;
      REGS_1909<=FA_cout_3444;
      REGS_1910<=FA_cout_3445;
      REGS_1911<=FA_cout_3446;
      REGS_1912<=FA_cout_3447;
      REGS_1913<=FA_cout_3448;
      REGS_1914<=FA_cout_3449;
      REGS_1915<=FA_cout_3450;
      REGS_1916<=FA_cout_3451;
      REGS_1917<=FA_cout_3452;
      REGS_1918<=FA_cout_3453;
      REGS_1919<=FA_cout_3454;
      REGS_1920<=FA_cout_3455;
      REGS_1921<=FA_cout_3456;
      REGS_1922<=FA_cout_3457;
      REGS_1923<=FA_cout_3458;
      REGS_1924<=FA_cout_3459;
      REGS_1925<=FA_cout_3460;
      REGS_1926<=FA_cout_3461;
      REGS_1927<=FA_cout_3462;
      REGS_1928<=FA_cout_3463;
      REGS_1929<=FA_cout_3464;
      REGS_1930<=FA_cout_3465;
      REGS_1931<=FA_cout_3466;
      REGS_1932<=FA_cout_3467;
      REGS_1933<=FA_cout_3468;
      REGS_1934<=FA_cout_3469;
      REGS_1935<=FA_cout_3470;
      REGS_1936<=FA_cout_3471;
      REGS_1937<=FA_cout_3472;
      REGS_1938<=FA_cout_3473;
      REGS_1939<=FA_cout_3474;
      REGS_1940<=FA_cout_3475;
      REGS_1941<=FA_cout_3476;
      REGS_1942<=FA_cout_3477;
      REGS_1943<=FA_cout_3478;
      REGS_1944<=FA_cout_3479;
      REGS_1945<=FA_cout_3480;
      REGS_1946<=FA_cout_3481;
      REGS_1947<=FA_cout_3482;
      REGS_1948<=FA_cout_3483;
      REGS_1949<=FA_cout_3484;
      REGS_1950<=FA_cout_3485;
      REGS_1951<=FA_cout_3486;
      REGS_1952<=FA_cout_3487;
      REGS_1953<=FA_cout_3488;
      REGS_1954<=FA_cout_3489;
      REGS_1955<=FA_cout_3490;
      REGS_1956<=FA_cout_3491;
      REGS_1957<=FA_cout_3492;
      REGS_1958<=FA_cout_3493;
      REGS_1959<=FA_cout_3494;
      REGS_1960<=FA_cout_3495;
      REGS_1961<=FA_cout_3496;
      REGS_1962<=FA_cout_3497;
      REGS_1963<=FA_cout_3498;
      REGS_1964<=HA_out_216;
      REGS_1965<=HA_out_217;
      REGS_1966<=HA_out_218;
      REGS_1967<=HA_out_219;
      REGS_1968<=HA_out_220;
      REGS_1969<=HA_out_221;
      REGS_1970<=HA_out_222;
      REGS_1971<=HA_out_223;
      REGS_1972<=FA_out_3444;
      REGS_1973<=FA_out_3445;
      REGS_1974<=FA_out_3446;
      REGS_1975<=FA_out_3447;
      REGS_1976<=FA_out_3448;
      REGS_1977<=FA_out_3449;
      REGS_1978<=FA_out_3450;
      REGS_1979<=FA_out_3451;
      REGS_1980<=FA_out_3452;
      REGS_1981<=FA_out_3453;
      REGS_1982<=FA_out_3454;
      REGS_1983<=FA_out_3455;
      REGS_1984<=FA_out_3456;
      REGS_1985<=FA_out_3457;
      REGS_1986<=FA_out_3458;
      REGS_1987<=FA_out_3459;
      REGS_1988<=FA_out_3460;
      REGS_1989<=FA_out_3461;
      REGS_1990<=FA_out_3462;
      REGS_1991<=FA_out_3463;
      REGS_1992<=FA_out_3464;
      REGS_1993<=FA_out_3465;
      REGS_1994<=FA_out_3466;
      REGS_1995<=FA_out_3467;
      REGS_1996<=FA_out_3468;
      REGS_1997<=FA_out_3469;
      REGS_1998<=FA_out_3470;
      REGS_1999<=FA_out_3471;
      REGS_2000<=FA_out_3472;
      REGS_2001<=FA_out_3473;
      REGS_2002<=FA_out_3474;
      REGS_2003<=FA_out_3475;
      REGS_2004<=FA_out_3476;
      REGS_2005<=FA_out_3477;
      REGS_2006<=FA_out_3478;
      REGS_2007<=FA_out_3479;
      REGS_2008<=FA_out_3480;
      REGS_2009<=FA_out_3481;
      REGS_2010<=FA_out_3482;
      REGS_2011<=FA_out_3483;
      REGS_2012<=FA_out_3484;
      REGS_2013<=FA_out_3485;
      REGS_2014<=FA_out_3486;
      REGS_2015<=FA_out_3487;
      REGS_2016<=FA_out_3488;
      REGS_2017<=FA_out_3489;
      REGS_2018<=FA_out_3490;
      REGS_2019<=FA_out_3491;
      REGS_2020<=FA_out_3492;
      REGS_2021<=FA_out_3493;
      REGS_2022<=FA_out_3494;
      REGS_2023<=FA_out_3495;
      REGS_2024<=FA_out_3496;
      REGS_2025<=FA_out_3497;
      REGS_2026<=FA_out_3498;
      REGS_2027<=FA_out_3499;
      REGS_2028<=FA_cout_3499;
      REGS_2029<=FA_out_3500;
      REGS_2030<=FA_cout_3500;
      REGS_2031<=FA_out_3501;
      REGS_2032<=FA_cout_3501;
      REGS_2033<=FA_out_3502;
      REGS_2034<=FA_cout_3502;
      REGS_2035<=FA_out_3503;
      REGS_2036<=FA_cout_3503;
      REGS_2037<=FA_out_3504;
      REGS_2038<=FA_cout_3504;
      REGS_2039<=HA_out_177;
      REGS_2040<=HA_out_178;
      REGS_2041<=HA_out_179;
      REGS_2042<=FA_out_3248;
      REGS_2043<=FA_out_3249;
      REGS_2044<=FA_out_3250;
      REGS_2045<=FA_out_3251;
      REGS_2046<=FA_out_3252;
      REGS_2047<=FA_out_3253;
      REGS_2048<=HA_out_224;
      REGS_2049<=HA_cout_224;
      REGS_2050<=HA_cout_225;
      REGS_2051<=HA_cout_226;
      REGS_2052<=HA_cout_227;
      REGS_2053<=FA_cout_3505;
      REGS_2054<=FA_cout_3506;
      REGS_2055<=FA_cout_3507;
      REGS_2056<=FA_cout_3508;
      REGS_2057<=FA_cout_3509;
      REGS_2058<=FA_cout_3510;
      REGS_2059<=FA_cout_3511;
      REGS_2060<=FA_cout_3512;
      REGS_2061<=FA_cout_3513;
      REGS_2062<=FA_cout_3514;
      REGS_2063<=FA_cout_3515;
      REGS_2064<=FA_cout_3516;
      REGS_2065<=FA_cout_3517;
      REGS_2066<=FA_cout_3518;
      REGS_2067<=FA_cout_3519;
      REGS_2068<=FA_cout_3520;
      REGS_2069<=FA_cout_3521;
      REGS_2070<=FA_cout_3522;
      REGS_2071<=FA_cout_3523;
      REGS_2072<=FA_cout_3524;
      REGS_2073<=FA_cout_3525;
      REGS_2074<=FA_cout_3526;
      REGS_2075<=FA_cout_3527;
      REGS_2076<=FA_cout_3528;
      REGS_2077<=FA_cout_3529;
      REGS_2078<=FA_cout_3530;
      REGS_2079<=FA_cout_3531;
      REGS_2080<=FA_cout_3532;
      REGS_2081<=FA_cout_3533;
      REGS_2082<=FA_cout_3534;
      REGS_2083<=FA_cout_3535;
      REGS_2084<=FA_cout_3536;
      REGS_2085<=FA_cout_3537;
      REGS_2086<=FA_cout_3538;
      REGS_2087<=FA_out_3539;
      REGS_2088<=FA_cout_3539;
      REGS_2089<=HA_out_225;
      REGS_2090<=HA_out_226;
      REGS_2091<=HA_out_227;
      REGS_2092<=FA_out_3505;
      REGS_2093<=FA_out_3506;
      REGS_2094<=FA_out_3507;
      REGS_2095<=FA_out_3508;
      REGS_2096<=FA_out_3509;
      REGS_2097<=FA_out_3510;
      REGS_2098<=FA_out_3511;
      REGS_2099<=FA_out_3512;
      REGS_2100<=FA_out_3513;
      REGS_2101<=FA_out_3514;
      REGS_2102<=FA_out_3515;
      REGS_2103<=FA_out_3516;
      REGS_2104<=FA_out_3517;
      REGS_2105<=FA_out_3518;
      REGS_2106<=FA_out_3519;
      REGS_2107<=FA_out_3520;
      REGS_2108<=FA_out_3521;
      REGS_2109<=FA_out_3522;
      REGS_2110<=FA_out_3523;
      REGS_2111<=FA_out_3524;
      REGS_2112<=FA_out_3525;
      REGS_2113<=FA_out_3526;
      REGS_2114<=FA_out_3527;
      REGS_2115<=FA_out_3528;
      REGS_2116<=FA_out_3529;
      REGS_2117<=FA_out_3530;
      REGS_2118<=FA_out_3531;
      REGS_2119<=FA_out_3532;
      REGS_2120<=FA_out_3533;
      REGS_2121<=FA_out_3534;
      REGS_2122<=FA_out_3535;
      REGS_2123<=FA_out_3536;
      REGS_2124<=FA_out_3537;
      REGS_2125<=FA_out_3538;
      REGS_2126<=FA_out_3540;
      REGS_2127<=FA_cout_3540;
      REGS_2128<=FA_out_3541;
      REGS_2129<=FA_cout_3541;
      REGS_2130<=FA_out_3542;
      REGS_2131<=FA_cout_3542;
      REGS_2132<=FA_out_3543;
      REGS_2133<=FA_cout_3543;
      REGS_2134<=FA_out_3544;
      REGS_2135<=FA_cout_3544;
      REGS_2136<=FA_out_3545;
      REGS_2137<=FA_cout_3545;
      REGS_2138<=FA_out_3546;
      REGS_2139<=FA_cout_3546;
      REGS_2140<=FA_out_3547;
      REGS_2141<=FA_cout_3547;
      REGS_2142<=FA_out_3548;
      REGS_2143<=FA_cout_3548;
      REGS_2144<=FA_out_3549;
      REGS_2145<=FA_cout_3549;
      REGS_2146<=FA_out_3550;
      REGS_2147<=FA_cout_3550;
      REGS_2148<=FA_out_3551;
      REGS_2149<=FA_cout_3551;
      REGS_2150<=FA_out_3552;
      REGS_2151<=FA_cout_3552;
      REGS_2152<=FA_out_3553;
      REGS_2153<=FA_cout_3553;
      REGS_2154<=FA_out_3554;
      REGS_2155<=FA_cout_3554;
      REGS_2156<=FA_out_3555;
      REGS_2157<=FA_cout_3555;
      REGS_2158<=FA_out_3556;
      REGS_2159<=FA_cout_3556;
      REGS_2160<=FA_out_3557;
      REGS_2161<=FA_cout_3557;
      REGS_2162<=FA_out_3558;
      REGS_2163<=FA_cout_3558;
      REGS_2164<=FA_out_3559;
      REGS_2165<=FA_cout_3559;
      REGS_2166<=FA_out_3560;
      REGS_2167<=FA_cout_3560;
      REGS_2168<=FA_out_3561;
      REGS_2169<=FA_cout_3561;
      REGS_2170<=FA_out_3562;
      REGS_2171<=FA_cout_3562;
      REGS_2172<=FA_out_3563;
      REGS_2173<=FA_cout_3563;
      REGS_2174<=FA_out_3564;
      REGS_2175<=FA_cout_3564;
      REGS_2176<=FA_out_3565;
      REGS_2177<=FA_cout_3565;
      REGS_2178<=FA_out_3566;
      REGS_2179<=FA_cout_3566;
      REGS_2180<=FA_out_3567;
      REGS_2181<=FA_cout_3567;
      REGS_2182<=FA_out_3568;
      REGS_2183<=FA_cout_3568;
      REGS_2184<=FA_out_3569;
      REGS_2185<=FA_cout_3569;
      REGS_2186<=FA_out_3570;
      REGS_2187<=FA_cout_3570;
      REGS_2188<=FA_out_3571;
      REGS_2189<=FA_cout_3571;
      REGS_2190<=FA_out_3572;
      REGS_2191<=FA_cout_3572;
      REGS_2192<=FA_out_3573;
      REGS_2193<=FA_cout_3573;
      REGS_2194<=FA_out_3574;
      REGS_2195<=FA_cout_3574;
      REGS_2196<=FA_out_3575;
      REGS_2197<=FA_cout_3575;
      REGS_2198<=FA_out_3576;
      REGS_2199<=FA_cout_3576;
      REGS_2200<=FA_out_3577;
      REGS_2201<=FA_cout_3577;
      REGS_2202<=FA_out_3578;
      REGS_2203<=FA_cout_3578;
      REGS_2204<=FA_out_3579;
      REGS_2205<=FA_cout_3579;
      REGS_2206<=FA_out_3580;
      REGS_2207<=FA_cout_3580;
      REGS_2208<=FA_out_3581;
      REGS_2209<=FA_cout_3581;
      REGS_2210<=FA_out_3582;
      REGS_2211<=FA_cout_3582;
      REGS_2212<=FA_out_3583;
      REGS_2213<=FA_cout_3583;
      REGS_2214<=FA_out_3584;
      REGS_2215<=FA_cout_3584;
      REGS_2216<=FA_out_3585;
      REGS_2217<=FA_cout_3585;
      REGS_2218<=FA_out_3586;
      REGS_2219<=FA_cout_3586;
      REGS_2220<=FA_out_3587;
      REGS_2221<=FA_cout_3587;
      REGS_2222<=FA_out_3588;
      REGS_2223<=FA_cout_3588;
      REGS_2224<=FA_out_3589;
      REGS_2225<=FA_cout_3589;
      REGS_2226<=FA_out_3590;
      REGS_2227<=FA_cout_3590;
      REGS_2228<=FA_out_3591;
      REGS_2229<=FA_cout_3591;
      REGS_2230<=FA_out_3592;
      REGS_2231<=FA_cout_3592;
      REGS_2232<=FA_out_3593;
      REGS_2233<=FA_cout_3593;
      REGS_2234<=FA_out_3594;
      REGS_2235<=FA_cout_3594;
      REGS_2236<=FA_out_3595;
      REGS_2237<=FA_cout_3595;
      REGS_2238<=HA_out_228;
      REGS_2239<=HA_cout_228;
      REGS_2240<=FA_out_3596;
      REGS_2241<=FA_cout_3596;
      REGS_2242<=HA_out_229;
      REGS_2243<=HA_cout_229;
      REGS_2244<=FA_out_3597;
      REGS_2245<=FA_cout_3597;
      REGS_2246<=HA_out_230;
      REGS_2247<=HA_cout_230;
      REGS_2248<=FA_out_3598;
      REGS_2249<=FA_cout_3598;
      REGS_2250<=HA_out_231;
      REGS_2251<=HA_cout_231;
      REGS_2252<=FA_out_3599;
      REGS_2253<=FA_cout_3599;
      REGS_2254<=HA_out_142;
      REGS_2255<=HA_out_143;
      REGS_2256<=HA_out_144;
      REGS_2257<=FA_out_3075;
      REGS_2258<=FA_out_3076;
      REGS_2259<=FA_out_3077;
      REGS_2260<=HA_out_187;
      REGS_2261<=HA_out_232;
      REGS_2262<=HA_cout_232;
      REGS_2263<=HA_cout_233;
      REGS_2264<=HA_cout_234;
      REGS_2265<=HA_cout_235;
      REGS_2266<=HA_cout_236;
      REGS_2267<=HA_cout_237;
      REGS_2268<=HA_cout_238;
      REGS_2269<=HA_cout_239;
      REGS_2270<=HA_cout_240;
      REGS_2271<=FA_cout_3600;
      REGS_2272<=FA_cout_3601;
      REGS_2273<=FA_cout_3602;
      REGS_2274<=FA_cout_3603;
      REGS_2275<=FA_cout_3604;
      REGS_2276<=FA_cout_3605;
      REGS_2277<=FA_cout_3606;
      REGS_2278<=HA_cout_241;
      REGS_2279<=FA_out_3411;
      REGS_2280<=FA_out_3607;
      REGS_2281<=FA_cout_3607;
      REGS_2282<=HA_out_233;
      REGS_2283<=HA_out_234;
      REGS_2284<=HA_out_235;
      REGS_2285<=HA_out_236;
      REGS_2286<=HA_out_237;
      REGS_2287<=HA_out_238;
      REGS_2288<=HA_out_239;
      REGS_2289<=HA_out_240;
      REGS_2290<=FA_out_3600;
      REGS_2291<=FA_out_3601;
      REGS_2292<=FA_out_3602;
      REGS_2293<=FA_out_3603;
      REGS_2294<=FA_out_3604;
      REGS_2295<=FA_out_3605;
      REGS_2296<=FA_out_3606;
      REGS_2297<=HA_out_241;
      REGS_2298<=HA_out_242;
      REGS_2299<=HA_cout_242;
      REGS_2300<=FA_out_3415;
      REGS_2301<=FA_out_3608;
      REGS_2302<=FA_cout_3608;
      REGS_2303<=HA_out_243;
      REGS_2304<=HA_cout_243;
      REGS_2305<=FA_out_3419;
      REGS_2306<=FA_out_3609;
      REGS_2307<=FA_cout_3609;
      REGS_2308<=HA_out_244;
      REGS_2309<=HA_cout_244;
      REGS_2310<=FA_out_3423;
      REGS_2311<=FA_out_3610;
      REGS_2312<=FA_cout_3610;
      REGS_2313<=HA_out_245;
      REGS_2314<=HA_cout_245;
      REGS_2315<=FA_out_3427;
      REGS_2316<=FA_out_3611;
      REGS_2317<=FA_cout_3611;
      REGS_2318<=HA_out_246;
      REGS_2319<=HA_cout_246;
      REGS_2320<=FA_out_3431;
      REGS_2321<=FA_out_3612;
      REGS_2322<=FA_cout_3612;
      REGS_2323<=HA_out_247;
      REGS_2324<=HA_cout_247;
      REGS_2325<=FA_out_3435;
      REGS_2326<=FA_out_3613;
      REGS_2327<=FA_cout_3613;
      REGS_2328<=HA_out_248;
      REGS_2329<=HA_cout_248;
      REGS_2330<=HA_out_191;
      REGS_2331<=HA_out_249;
      REGS_2332<=HA_cout_249;
      REGS_2333<=HA_out_250;
      REGS_2334<=HA_cout_250;
      REGS_2335<=FA_out_3152;
      REGS_2336<=HA_out_251;
      REGS_2337<=HA_cout_251;
      REGS_2338<=HA_out_252;
      REGS_2339<=HA_cout_252;
      REGS_2340<=HA_out_253;
      REGS_2341<=HA_cout_253;
      REGS_2342<=HA_out_254;
      REGS_2343<=HA_cout_254;
      REGS_2344<=HA_out_255;
      REGS_2345<=HA_cout_255;
      REGS_2346<=HA_out_256;
      REGS_2347<=HA_cout_256;
      REGS_2348<=HA_out_257;
      REGS_2349<=HA_cout_257;
      REGS_2350<=HA_out_258;
      REGS_2351<=HA_cout_258;
      REGS_2352<=HA_out_259;
      REGS_2353<=HA_cout_259;
      REGS_2354<=HA_out_260;
      REGS_2355<=HA_cout_260;
      REGS_2356<=FA_out_3182;
      REGS_2357<=HA_out_261;
      REGS_2358<=HA_cout_261;
      REGS_2359<=HA_out_153;
      REGS_2360<=HA_out_262;
      REGS_2361<=HA_cout_262;
      REGS_2362<=HA_out_157;
      REGS_2363<=HA_out_263;
      REGS_2364<=HA_cout_263;
      REGS_2365<=HA_out_160;
      REGS_2366<=HA_out_264;
      REGS_2367<=HA_cout_264;
      REGS_2368<=HA_out_165;
      REGS_2369<=HA_out_265;
      REGS_2370<=HA_cout_265;
      REGS_2371<=HA_out_212;
      REGS_2372<=HA_out_168;
      REGS_2373<=HA_out_266;
      REGS_2374<=HA_cout_266;
      REGS_2375<=REGS_1842;
      REGS_2376<=REGS_1888;
  end


endmodule

